configuration coin_register_behaviour_cfg of coin_register is
   for behaviour
   end for;
end coin_register_behaviour_cfg;

library IEEE;
use IEEE.std_logic_1164.ALL;

entity video_system_tb is
end video_system_tb;


configuration shift_ctrl_gg_behaviour_cfg of shift_ctrl_gg is
   for behaviour
   end for;
end shift_ctrl_gg_behaviour_cfg;

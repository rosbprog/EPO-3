library IEEE;
use IEEE.std_logic_1164.ALL;

entity ghost_cont_tb is
end ghost_cont_tb;


configuration coordinate_register_behavioural_cfg of coordinate_register is
   for behavioural
   end for;
end coordinate_register_behavioural_cfg;

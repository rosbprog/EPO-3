configuration shift_ctrl_gr_behaviour_cfg of shift_ctrl_gr is
   for behaviour
   end for;
end shift_ctrl_gr_behaviour_cfg;

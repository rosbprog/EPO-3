configuration multiplexer_behaviour_cfg of multiplexer is
   for behaviour
   end for;
end multiplexer_behaviour_cfg;

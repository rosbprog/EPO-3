configuration coordinate_adder_behavioural_cfg of coordinate_adder is
   for behavioural
   end for;
end coordinate_adder_behavioural_cfg;

configuration shift_counter_behaviour_cfg of shift_counter is
   for behaviour
   end for;
end shift_counter_behaviour_cfg;

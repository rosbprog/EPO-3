configuration video_counter_behaviour_cfg of video_counter is
   for behaviour
   end for;
end video_counter_behaviour_cfg;

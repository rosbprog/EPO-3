configuration cell_register_behavioural_cfg of cell_register is
   for behavioural
   end for;
end cell_register_behavioural_cfg;

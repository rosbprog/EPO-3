library IEEE;
use IEEE.std_logic_1164.ALL;

entity shift_system_tb is
end shift_system_tb;


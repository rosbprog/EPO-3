configuration counter_behavioural_cfg of counter is
   for behavioural
   end for;
end counter_behavioural_cfg;

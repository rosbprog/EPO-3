configuration vga_controll_vga_behavioral_cfg of vga_controll is
   for vga_behavioral
   end for;
end vga_controll_vga_behavioral_cfg;

configuration gr_pos_reg_behaviour_cfg of gr_pos_reg is
   for behaviour
   end for;
end gr_pos_reg_behaviour_cfg;

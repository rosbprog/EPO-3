configuration shift_count_gg_behaviour_cfg of shift_count_gg is
   for behaviour
   end for;
end shift_count_gg_behaviour_cfg;

configuration coordinate_comparator_behavioural_cfg of coordinate_comparator is
   for behavioural
   end for;
end coordinate_comparator_behavioural_cfg;

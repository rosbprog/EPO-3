configuration fsm_counter_behavioural_cfg of fsm_counter is
   for behavioural
   end for;
end fsm_counter_behavioural_cfg;

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity pacman_position_reg_tb is
end entity;

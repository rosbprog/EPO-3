configuration gameover_control_behaviour_cfg of gameover_control is
   for behaviour
   end for;
end gameover_control_behaviour_cfg;

configuration score_count_behaviour_cfg of score_count is
   for behaviour
   end for;
end score_count_behaviour_cfg;

configuration pulse_generator_behavioural_cfg of pulse_generator is
   for behavioural
   end for;
end pulse_generator_behavioural_cfg;

library IEEE;
use IEEE.std_logic_1164.all;

entity buffer_1bit is
	port (	
		clk	:in  std_logic;
		input	:in  std_logic;
		output	:out std_logic
	);
end entity buffer_1bit;	



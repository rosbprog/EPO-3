library IEEE;
use IEEE.std_logic_1164.all;

entity sprite is
	port(  	y_pos		:in std_logic_vector (2 downto 0); 
		--Upper row is 111, lower is 000
	 	sprite_select	:in std_logic_vector (2 downto 0); 
		--000 coin, 001 ghost_red, 010 ghost_green, 011 pacman, 100 wall
		--What do we chose when accidentally e.g. 101 gets sampled? now pacman.
		color_out 	:out std_logic_vector (2 downto 0); --respectively RGB	
		row_out		:out std_logic_vector (7 downto 0)  --left to right		
		);
end entity sprite;

architecture behavioural of sprite is
begin
	process(y_pos, sprite_select)
		begin
			if(sprite_select = "000") then  --coin
				color_out <= "111";
				if(y_pos = "111") then
					row_out <= "00000000"; 
				elsif(y_pos = "110") then
					row_out <= "00000000"; 
				elsif(y_pos = "101") then
					row_out <= "00011000";
				elsif(y_pos = "100") then
					row_out <= "00111100";
				elsif(y_pos = "011") then
					row_out <= "00111100";
				elsif(y_pos = "010") then
					row_out <= "00011000";
				elsif(y_pos = "001") then
					row_out <= "00000000";
				else
					row_out <= "00000000";
				end if; 
			
			elsif(sprite_select = "001") then  --wall
				color_out <= "001";
				if(y_pos = "111") then
					row_out <= "11111111"; 
				elsif(y_pos = "110") then
					row_out <= "11111111"; 
				elsif(y_pos = "101") then
					row_out <= "11111111";
				elsif(y_pos = "100") then
					row_out <= "11111111";
				elsif(y_pos = "011") then
					row_out <= "11111111";
				elsif(y_pos = "010") then
					row_out <= "11111111";
				elsif(y_pos = "001") then
					row_out <= "11111111";
				else
					row_out <= "11111111";
				end if; 
			
			elsif(sprite_select = "010") then  --ghost red
				color_out <= "100";
				if(y_pos = "111") then
					row_out <= "00000000"; 
				elsif(y_pos = "110") then
					row_out <= "00111100"; 
				elsif(y_pos = "101") then
					row_out <= "01111110";
				elsif(y_pos = "100") then
					row_out <= "01011010";
				elsif(y_pos = "011") then
					row_out <= "01111110";
				elsif(y_pos = "010") then
					row_out <= "01111110";
				elsif(y_pos = "001") then
					row_out <= "01011010";
				else
					row_out <= "00000000";
				end if; 

			elsif(sprite_select = "011") then  --ghost green
				color_out <= "010";
				if(y_pos = "111") then
					row_out <= "00000000"; 
				elsif(y_pos = "110") then
					row_out <= "00111100"; 
				elsif(y_pos = "101") then
					row_out <= "01111110";
				elsif(y_pos = "100") then
					row_out <= "01011010";
				elsif(y_pos = "011") then
					row_out <= "01111110";
				elsif(y_pos = "010") then
					row_out <= "01111110";
				elsif(y_pos = "001") then
					row_out <= "01011010";
				else
					row_out <= "00000000";
				end if; 

			else  				--pacman
				color_out <= "110";
				if(y_pos = "111") then
					row_out <= "00000000"; 
				elsif(y_pos = "110") then
					row_out <= "00111100"; 
				elsif(y_pos = "101") then
					row_out <= "01110110";
				elsif(y_pos = "100") then
					row_out <= "01111110";
				elsif(y_pos = "011") then
					row_out <= "01111000";
				elsif(y_pos = "010") then
					row_out <= "01111110";
				elsif(y_pos = "001") then
					row_out <= "00111100";
				else
					row_out <= "00000000";
				end if;
			end if; 
	end process;
end architecture behavioural;


					
				
				
					

				


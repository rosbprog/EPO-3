configuration gg_pos_reg_behaviour_cfg of gg_pos_reg is
   for behaviour
   end for;
end gg_pos_reg_behaviour_cfg;

configuration row_controller_behavioural_cfg of row_controller is
   for behavioural
   end for;
end row_controller_behavioural_cfg;

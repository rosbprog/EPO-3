configuration ghost_cont_behaviour_cfg of ghost_cont is
   for behaviour
   end for;
end ghost_cont_behaviour_cfg;

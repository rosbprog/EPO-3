configuration vga_controll_tb_behaviour_cfg of vga_controll_tb is
   for behaviour
      for all: vga_controll use configuration work.vga_controll_vga_behavioral_cfg;
      end for;
   end for;
end vga_controll_tb_behaviour_cfg;

configuration video_control_behaviour_cfg of video_control is
   for behaviour
   end for;
end video_control_behaviour_cfg;

configuration shift_count_gr_behaviour_cfg of shift_count_gr is
   for behaviour
   end for;
end shift_count_gr_behaviour_cfg;

configuration reset_controller_behavioural_cfg of reset_controller is
   for behavioural
   end for;
end reset_controller_behavioural_cfg;

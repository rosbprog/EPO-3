configuration game_struct_tb_structural_cfg of game_struct_tb is
   for structural
      for all: game_struct use configuration work.game_struct_structural_cfg;
      end for;
   end for;
end game_struct_tb_structural_cfg;

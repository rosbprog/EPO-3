configuration score_control_behaviour_cfg of score_control is
   for behaviour
   end for;
end score_control_behaviour_cfg;

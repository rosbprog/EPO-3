configuration screen_controller_behavioural_cfg of screen_controller is
   for behavioural
   end for;
end screen_controller_behavioural_cfg;

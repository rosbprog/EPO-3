library IEEE;
use IEEE.std_logic_1164.ALL;

entity video_c_c_tb is
end video_c_c_tb;


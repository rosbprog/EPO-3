library IEEE;
use IEEE.std_logic_1164.ALL;

entity vc_tb is
end vc_tb;


library IEEE;
use IEEE.std_logic_1164.ALL;

entity score_counter_tb is
end score_counter_tb;


configuration counter_behaviour_cfg of counter is
   for behaviour
   end for;
end counter_behaviour_cfg;

configuration character_sprite_behavioural_cfg of character_sprite is
   for behavioural
   end for;
end character_sprite_behavioural_cfg;

configuration d_flip_flop_behavioural_cfg of d_flip_flop is
   for behavioural
   end for;
end d_flip_flop_behavioural_cfg;

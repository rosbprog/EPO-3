configuration sprite_behaviour_cfg of sprite is
   for behaviour
   end for;
end sprite_behaviour_cfg;

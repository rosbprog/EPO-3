configuration sprites_behaviour_cfg of sprites is
   for behaviour
   end for;
end sprites_behaviour_cfg;

configuration input_controller_behavioural_cfg of input_controller is
   for behavioural
   end for;
end input_controller_behavioural_cfg;

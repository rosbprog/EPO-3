configuration coordinate_multiplexer_behavioural_cfg of coordinate_multiplexer is
   for behavioural
   end for;
end coordinate_multiplexer_behavioural_cfg;

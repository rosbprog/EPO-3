configuration map_register_behaviour_cfg of map_register is
   for behaviour
      for all: row_controller use configuration work.row_controller_behavioural_cfg;
      end for;
   end for;
end map_register_behaviour_cfg;

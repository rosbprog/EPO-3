library IEEE;
use IEEE.std_logic_1164.ALL;

entity vga_controll_tb is
end vga_controll_tb;



library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of total_system is

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AO31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component EDFKCND1BWP7T
    port(CP, CN, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component OA222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component EDFKCNQD1BWP7T
    port(CP, CN, D, E : in std_logic; Q : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component DFXD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKCND0BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component BUFFD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DFQD0BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component MUX2D0BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component DFKSND1BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AO33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component MUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component OR4XD1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component OR3XD1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component NR3D1BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component LNQD1BWP7T
    port(EN, D : in std_logic; Q : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  signal cell_type_int : std_logic_vector(2 downto 0);
  signal L1_row_new_pacman : std_logic_vector(4 downto 0);
  signal ycoordinates_int : std_logic_vector(4 downto 0);
  signal L1_row_old_ghost1 : std_logic_vector(4 downto 0);
  signal L1_col_new_pacman : std_logic_vector(4 downto 0);
  signal xcoordinates_int : std_logic_vector(4 downto 0);
  signal L1_col_old_ghost1 : std_logic_vector(4 downto 0);
  signal L1_L3a_move : std_logic_vector(3 downto 0);
  signal L1_row_old_pacman : std_logic_vector(4 downto 0);
  signal L1_col_old_pacman : std_logic_vector(4 downto 0);
  signal L1_L3a_L5_state : std_logic_vector(1 downto 0);
  signal L1_L1a_coin_memory : std_logic_vector(47 downto 0);
  signal L1_row_coin : std_logic_vector(4 downto 0);
  signal L1_col_coin : std_logic_vector(4 downto 0);
  signal L1_L3b_L5_state : std_logic_vector(1 downto 0);
  signal L1_L3c_move : std_logic_vector(3 downto 0);
  signal L1_L3c_PC1_state : std_logic_vector(2 downto 0);
  signal L1_L6a_LBL1_state : std_logic_vector(3 downto 0);
  signal L1_L6a_LBL2_count : std_logic_vector(6 downto 0);
  signal L1_L3a_L0_data_intermediate : std_logic_vector(3 downto 0);
  signal L1_L3a_data_buffed : std_logic_vector(3 downto 0);
  signal L2_vgacontrol_hcount : std_logic_vector(9 downto 0);
  signal L2_vgacontrol_vcount : std_logic_vector(9 downto 0);
  signal L2_screencontrol_state : std_logic_vector(1 downto 0);
  signal L2_in_go_sprite_type : std_logic_vector(4 downto 0);
  signal L2_in_go_colour : std_logic_vector(2 downto 0);
  signal L2_rgb_score : std_logic_vector(2 downto 0);
  signal L2_rgb_video : std_logic_vector(2 downto 0);
  signal L2_score_score_sprite_type : std_logic_vector(3 downto 0);
  signal L2_in_go_y_pos : std_logic_vector(2 downto 0);
  signal L2_county : std_logic_vector(2 downto 0);
  signal L2_shift_L12_count_internal : std_logic_vector(2 downto 0);
  signal L2_shift_pixel_arr_out_shift_gg : std_logic_vector(7 downto 0);
  signal L2_shift_pixel_arr_out_shift_gr : std_logic_vector(7 downto 0);
  signal L2_shift_pixel_arr_out_shift_pacman : std_logic_vector(7 downto 0);
  signal L2_pixel_array_shifted : std_logic_vector(7 downto 0);
  signal L2_pixel_array_to_shift : std_logic_vector(7 downto 0);
  signal L2_shift_cell_state_out_shift_pacman : std_logic_vector(5 downto 0);
  signal L2_sprite_colour : std_logic_vector(2 downto 0);
  signal L2_shift_y_pos_out_shift_pacman : std_logic_vector(2 downto 0);
  signal L2_shift_y_pos_out_shift_gg : std_logic_vector(2 downto 0);
  signal L2_shift_y_pos_out_shift_gr : std_logic_vector(2 downto 0);
  signal L2_shift_cell_state_out_shift_gr : std_logic_vector(2 downto 0);
  signal L2_shift_cell_state_out_shift_gg : std_logic_vector(2 downto 0);
  signal L2_current_block_horizontal : std_logic_vector(4 downto 0);
  signal L2_current_block_vertical : std_logic_vector(4 downto 0);
  signal L2_shift_pacman_pos_x : std_logic_vector(4 downto 0);
  signal L2_shift_pacman_pos_y : std_logic_vector(4 downto 0);
  signal L2_shift_gr_pos_x : std_logic_vector(4 downto 0);
  signal L2_shift_gr_pos_y : std_logic_vector(4 downto 0);
  signal L2_shift_gg_pos_x : std_logic_vector(4 downto 0);
  signal L2_shift_gg_pos_y : std_logic_vector(4 downto 0);
  signal L2_shift_pacman_pos_x_new : std_logic_vector(4 downto 0);
  signal L2_shift_gr_pos_x_new : std_logic_vector(4 downto 0);
  signal L2_shift_pacman_pos_y_new : std_logic_vector(4 downto 0);
  signal L2_shift_gr_pos_y_new : std_logic_vector(4 downto 0);
  signal L2_shift_gg_pos_x_new : std_logic_vector(4 downto 0);
  signal L2_shift_gg_pos_y_new : std_logic_vector(4 downto 0);
  signal L2_shift_L31_count_internal : std_logic_vector(2 downto 0);
  signal L2_shift_L33_state : std_logic_vector(4 downto 0);
  signal L2_shift_L21_count_internal : std_logic_vector(2 downto 0);
  signal L2_shift_L23_state : std_logic_vector(4 downto 0);
  signal L2_in_score_12bits : std_logic_vector(11 downto 0);
  signal L2_gameovercontrol_state : std_logic_vector(3 downto 0);
  signal L2_gameovercontrol_pixel_arr_buffer : std_logic_vector(7 downto 0);
  signal L2_score_L3_pixel_arr_buffer : std_logic_vector(7 downto 0);
  signal L2_score_L3_state : std_logic_vector(3 downto 0);
  signal L2_shift_L11_state : std_logic_vector(4 downto 0);
  signal L1_L6b_state : std_logic_vector(1 downto 0);
  signal L1_L3c_IS1_IC1_state : std_logic_vector(2 downto 0);
  signal L1_L3c_IS1_data_intermediate : std_logic_vector(3 downto 0);
  signal L1_L3a_L1_state : std_logic_vector(2 downto 0);
  signal L2_vidcontrol_colour_buffer : std_logic_vector(2 downto 0);
  signal L2_vidcontrol_pixel_arr_buffer : std_logic_vector(7 downto 0);
  signal L2_vidcontrol_state : std_logic_vector(3 downto 0);
  signal L1_L3c_IS1_IB1_data_intermediate : std_logic_vector(3 downto 0);
  signal L1_L1a_n_0, L1_L1a_n_1, L1_L1a_n_2, L1_L1a_n_3, L1_L1a_n_5 : std_logic;
  signal L1_L1a_n_6, L1_L1a_n_7, L1_L1a_n_8, L1_L1a_n_9, L1_L1a_n_10 : std_logic;
  signal L1_L1a_n_11, L1_L1a_n_12, L1_L1a_n_13, L1_L1a_n_14, L1_L1a_n_16 : std_logic;
  signal L1_L1a_n_17, L1_L1a_n_18, L1_L1a_n_19, L1_L1a_n_20, L1_L1a_n_21 : std_logic;
  signal L1_L1a_n_22, L1_L1a_n_23, L1_L1a_n_24, L1_L1a_n_25, L1_L1a_n_26 : std_logic;
  signal L1_L1a_n_27, L1_L1a_n_28, L1_L1a_n_29, L1_L1a_n_30, L1_L1a_n_31 : std_logic;
  signal L1_L1a_n_32, L1_L1a_n_33, L1_L1a_n_34, L1_L1a_n_35, L1_L1a_n_36 : std_logic;
  signal L1_L1a_n_37, L1_L1a_n_38, L1_L1a_n_39, L1_L1a_n_40, L1_L1a_n_41 : std_logic;
  signal L1_L1a_n_42, L1_L1a_n_43, L1_L1a_n_44, L1_L1a_n_45, L1_L1a_n_46 : std_logic;
  signal L1_L1a_n_47, L1_L1a_n_48, L1_L1a_n_49, L1_L1a_n_50, L1_L1a_n_51 : std_logic;
  signal L1_L1a_n_52, L1_L1a_n_53, L1_L1a_n_54, L1_L1a_n_55, L1_L1a_n_56 : std_logic;
  signal L1_L1a_n_57, L1_L1a_n_58, L1_L1a_n_59, L1_L1a_n_60, L1_L1a_n_61 : std_logic;
  signal L1_L1a_n_62, L1_L1a_n_63, L1_L1a_n_64, L1_L1a_n_65, L1_L1a_n_66 : std_logic;
  signal L1_L1a_n_67, L1_L1a_n_68, L1_L1a_n_69, L1_L1a_n_70, L1_L1a_n_71 : std_logic;
  signal L1_L1a_n_72, L1_L1a_n_73, L1_L1a_n_74, L1_L1a_n_75, L1_L1a_n_76 : std_logic;
  signal L1_L1a_n_77, L1_L1a_n_78, L1_L1a_n_79, L1_L1a_n_80, L1_L1a_n_81 : std_logic;
  signal L1_L1a_n_82, L1_L1a_n_83, L1_L1a_n_84, L1_L1a_n_85, L1_L1a_n_86 : std_logic;
  signal L1_L1a_n_87, L1_L1a_n_88, L1_L1a_n_89, L1_L1a_n_90, L1_L1a_n_91 : std_logic;
  signal L1_L1a_n_92, L1_L1a_n_93, L1_L1a_n_94, L1_L1a_n_95, L1_L1a_n_96 : std_logic;
  signal L1_L1a_n_97, L1_L1a_n_98, L1_L1a_n_99, L1_L1a_n_100, L1_L1a_n_101 : std_logic;
  signal L1_L1a_n_102, L1_L1a_n_103, L1_L1a_n_104, L1_L1a_n_105, L1_L1a_n_106 : std_logic;
  signal L1_L1a_n_107, L1_L1a_n_108, L1_L1a_n_109, L1_L1a_n_110, L1_L1a_n_111 : std_logic;
  signal L1_L1a_n_112, L1_L1a_n_113, L1_L1a_n_114, L1_L1a_n_115, L1_L1a_n_116 : std_logic;
  signal L1_L1a_n_117, L1_L1a_n_118, L1_L1a_n_119, L1_L1a_n_120, L1_L1a_n_121 : std_logic;
  signal L1_L1a_n_122, L1_L1a_n_123, L1_L1a_n_124, L1_L1a_n_125, L1_L1a_n_126 : std_logic;
  signal L1_L1a_n_127, L1_L1a_n_128, L1_L1a_n_129, L1_L1a_n_130, L1_L1a_n_131 : std_logic;
  signal L1_L1a_n_132, L1_L1a_n_133, L1_L1a_n_134, L1_L1a_n_135, L1_L1a_n_136 : std_logic;
  signal L1_L1a_n_137, L1_L1a_n_138, L1_L1a_n_139, L1_L1a_n_140, L1_L1a_n_141 : std_logic;
  signal L1_L1a_n_142, L1_L1a_n_143, L1_L1a_n_144, L1_L1a_n_145, L1_L1a_n_146 : std_logic;
  signal L1_L1a_n_147, L1_L1a_n_148, L1_L1a_n_149, L1_L1a_n_150, L1_L1a_n_151 : std_logic;
  signal L1_L1a_n_152, L1_L1a_n_153, L1_L1a_n_154, L1_L1a_n_155, L1_L1a_n_156 : std_logic;
  signal L1_L1a_n_157, L1_L1a_n_158, L1_L1a_n_159, L1_L1a_n_160, L1_L1a_n_161 : std_logic;
  signal L1_L1a_n_162, L1_L1a_n_163, L1_L1a_n_164, L1_L1a_n_165, L1_L1a_n_166 : std_logic;
  signal L1_L1a_n_167, L1_L1a_n_168, L1_L1a_n_169, L1_L1a_n_170, L1_L1a_n_171 : std_logic;
  signal L1_L1a_n_172, L1_L1a_n_173, L1_L1a_n_174, L1_L1a_n_175, L1_L1a_n_176 : std_logic;
  signal L1_L1a_n_177, L1_L1a_n_178, L1_L1a_n_179, L1_L1a_n_180, L1_L1a_n_181 : std_logic;
  signal L1_L1a_n_182, L1_L1a_n_183, L1_L1a_n_184, L1_L1a_n_185, L1_L1a_n_186 : std_logic;
  signal L1_L1a_n_187, L1_L1a_n_188, L1_L1a_n_189, L1_L1a_n_190, L1_L1a_n_191 : std_logic;
  signal L1_L1a_n_192, L1_L1a_n_193, L1_L1a_n_194, L1_L1a_n_195, L1_L1a_n_196 : std_logic;
  signal L1_L1a_n_197, L1_L1a_n_198, L1_L1a_n_199, L1_L1a_n_200, L1_L1a_n_201 : std_logic;
  signal L1_L1a_n_202, L1_L1a_n_203, L1_L1a_n_204, L1_L1a_n_206, L1_L1a_n_224 : std_logic;
  signal L1_L1a_n_225, L1_L1b_n_0, L1_L2_IB1_n_0, L1_L2_IB1_n_1, L1_L2_IB1_n_2 : std_logic;
  signal L1_L2_IB1_n_3, L1_L2_IB1_n_4, L1_L2_IB1_n_5, L1_L2_IB1_n_6, L1_L2_IB1_n_7 : std_logic;
  signal L1_L2_IB1_n_8, L1_L2_IB1_n_9, L1_L2_IB1_n_10, L1_L2_IB1_n_11, L1_L2_IB2_n_0 : std_logic;
  signal L1_L2_IB2_n_1, L1_L2_c_g1, L1_L2_c_g2, L1_L3a_L0_FF1_n_0, L1_L3a_L0_FF2_n_0 : std_logic;
  signal L1_L3a_L1_n_1, L1_L3a_L1_n_3, L1_L3a_L1_n_4, L1_L3a_L1_n_5, L1_L3a_L1_n_7 : std_logic;
  signal L1_L3a_L1_n_9, L1_L3a_L1_n_10, L1_L3a_L1_n_12, L1_L3a_L1_n_13, L1_L3a_L1_n_14 : std_logic;
  signal L1_L3a_L1_n_15, L1_L3a_L1_n_16, L1_L3a_L1_n_17, L1_L3a_L1_n_19, L1_L3a_L1_n_20 : std_logic;
  signal L1_L3a_L1_n_21, L1_L3a_L1_n_22, L1_L3a_L1_n_23, L1_L3a_L1_n_24, L1_L3a_L1_n_25 : std_logic;
  signal L1_L3a_L1_n_26, L1_L3a_L1_n_27, L1_L3a_L1_n_34, L1_L3a_L1_n_35, L1_L3a_L1_n_36 : std_logic;
  signal L1_L3a_L1_n_37, L1_L3a_L1_n_38, L1_L3b_n_0, L1_L3b_n_1, L1_L3b_n_2 : std_logic;
  signal L1_L3b_n_5, L1_L3b_n_6, L1_L3c_IS1_IB1_FF1_n_0, L1_L3c_IS1_IB1_FF2_n_0, L1_L3c_IS1_IC1_n_1 : std_logic;
  signal L1_L3c_IS1_IC1_n_2, L1_L3c_IS1_IC1_n_3, L1_L3c_IS1_IC1_n_4, L1_L3c_IS1_IC1_n_5, L1_L3c_IS1_IC1_n_6 : std_logic;
  signal L1_L3c_IS1_IC1_n_7, L1_L3c_IS1_IC1_n_8, L1_L3c_IS1_IC1_n_9, L1_L3c_IS1_IC1_n_11, L1_L3c_IS1_IC1_n_12 : std_logic;
  signal L1_L3c_IS1_IC1_n_15, L1_L3c_IS1_IC1_n_16, L1_L3c_IS1_IC1_n_17, L1_L3c_IS1_IC1_n_18, L1_L3c_IS1_IC1_n_19 : std_logic;
  signal L1_L3c_IS1_IC1_n_20, L1_L3c_IS1_IC1_n_21, L1_L3c_IS1_IC1_n_22, L1_L3c_IS1_IC1_n_23, L1_L3c_IS1_IC1_n_24 : std_logic;
  signal L1_L3c_IS1_IC1_n_25, L1_L3c_IS1_IC1_n_26, L1_L3c_IS1_IC1_n_27, L1_L3c_IS1_IC1_n_34, L1_L3c_IS1_IC1_n_36 : std_logic;
  signal L1_L3c_PC1_n_0, L1_L3c_PC1_n_1, L1_L3c_PC1_n_2, L1_L3c_PC1_n_3, L1_L3c_PC1_n_4 : std_logic;
  signal L1_L3c_PC1_n_5, L1_L3c_PC1_n_7, L1_L3c_PC1_n_8, L1_L3c_PC1_n_9, L1_L3c_n_0 : std_logic;
  signal L1_L3c_n_1, L1_L3c_n_2, L1_L3c_n_3, L1_L3c_n_4, L1_L3c_n_5 : std_logic;
  signal L1_L3c_n_6, L1_L3c_n_7, L1_L3c_n_8, L1_L3c_n_9, L1_L3c_n_10 : std_logic;
  signal L1_L3c_n_11, L1_L3c_n_12, L1_L3c_n_13, L1_L3c_n_14, L1_L3c_n_15 : std_logic;
  signal L1_L3c_n_16, L1_L3c_n_17, L1_L3c_n_18, L1_L3c_n_19, L1_L3c_n_20 : std_logic;
  signal L1_L3c_n_21, L1_L3c_n_22, L1_L3c_n_23, L1_L3c_n_24, L1_L3c_n_25 : std_logic;
  signal L1_L3c_n_26, L1_L3c_n_27, L1_L3c_n_28, L1_L3c_n_29, L1_L3c_n_30 : std_logic;
  signal L1_L3c_n_31, L1_L3c_n_32, L1_L3c_n_33, L1_L3c_n_34, L1_L3c_n_35 : std_logic;
  signal L1_L3c_n_36, L1_L3c_n_37, L1_L3c_n_38, L1_L3c_n_39, L1_L3c_n_40 : std_logic;
  signal L1_L3c_n_41, L1_L3c_n_42, L1_L3c_n_43, L1_L3c_n_44, L1_L3c_n_45 : std_logic;
  signal L1_L3c_n_46, L1_L3c_n_47, L1_L3c_n_48, L1_L3c_n_49, L1_L3c_n_50 : std_logic;
  signal L1_L3c_n_51, L1_L3c_n_52, L1_L3c_n_53, L1_L3c_n_54, L1_L3c_n_55 : std_logic;
  signal L1_L3c_n_56, L1_L3c_n_57, L1_L3c_n_58, L1_L3c_n_59, L1_L3c_n_60 : std_logic;
  signal L1_L3c_n_61, L1_L5_n_14, L1_L6a_LBL1_n_2, L1_L6a_LBL1_n_3, L1_L6a_LBL1_n_4 : std_logic;
  signal L1_L6a_LBL1_n_5, L1_L6a_LBL1_n_6, L1_L6a_LBL1_n_7, L1_L6a_LBL1_n_8, L1_L6a_LBL1_n_9 : std_logic;
  signal L1_L6a_LBL1_n_10, L1_L6a_LBL1_n_11, L1_L6a_LBL1_n_12, L1_L6a_LBL1_n_14, L1_L6a_LBL1_n_15 : std_logic;
  signal L1_L6a_LBL1_n_16, L1_L6a_LBL1_n_17, L1_L6a_LBL1_n_18, L1_L6a_LBL1_n_19, L1_L6a_LBL1_n_20 : std_logic;
  signal L1_L6a_LBL1_n_21, L1_L6a_LBL1_n_22, L1_L6a_LBL1_n_23, L1_L6a_LBL1_n_24, L1_L6a_LBL1_n_25 : std_logic;
  signal L1_L6a_LBL1_n_26, L1_L6a_LBL1_n_27, L1_L6a_LBL1_n_29, L1_L6a_LBL1_n_30, L1_L6a_LBL1_n_31 : std_logic;
  signal L1_L6a_LBL1_n_32, L1_L6a_LBL1_n_33, L1_L6a_LBL1_n_34, L1_L6a_LBL1_n_35, L1_L6a_LBL1_n_36 : std_logic;
  signal L1_L6a_LBL1_n_38, L1_L6a_LBL1_n_39, L1_L6a_LBL1_n_40, L1_L6a_LBL1_n_41, L1_L6a_LBL1_n_42 : std_logic;
  signal L1_L6a_LBL1_n_43, L1_L6a_LBL1_n_44, L1_L6a_LBL1_n_45, L1_L6a_LBL1_n_46, L1_L6a_LBL1_n_47 : std_logic;
  signal L1_L6a_LBL1_n_48, L1_L6a_LBL1_n_49, L1_L6a_LBL1_n_50, L1_L6a_LBL1_n_51, L1_L6a_LBL1_n_52 : std_logic;
  signal L1_L6a_LBL1_n_53, L1_L6a_LBL1_n_54, L1_L6a_LBL1_n_55, L1_L6a_LBL1_n_56, L1_L6a_LBL1_n_57 : std_logic;
  signal L1_L6a_LBL1_n_62, L1_L6a_LBL1_n_63, L1_L6a_LBL1_n_64, L1_L6a_LBL1_n_65, L1_L6a_LBL1_n_74 : std_logic;
  signal L1_L6a_LBL1_n_75, L1_L6a_LBL1_n_76, L1_L6a_LBL2_n_0, L1_L6a_LBL2_n_1, L1_L6a_LBL2_n_2 : std_logic;
  signal L1_L6a_LBL2_n_3, L1_L6a_LBL2_n_4, L1_L6a_LBL2_n_6, L1_L6a_LBL2_n_7, L1_L6a_LBL2_n_8 : std_logic;
  signal L1_L6a_LBL2_n_9, L1_L6a_LBL2_n_10, L1_L6a_LBL2_n_11, L1_L6a_LBL2_n_12, L1_L6a_LBL2_n_13 : std_logic;
  signal L1_L6a_LBL2_n_14, L1_L6a_LBL2_n_15, L1_L6a_LBL2_n_16, L1_L6a_LBL2_n_17, L1_L6a_LBL2_n_18 : std_logic;
  signal L1_L6a_LBL2_n_19, L1_L6a_LBL2_n_20, L1_L6a_LBL2_n_21, L1_L6a_LBL2_n_22, L1_L6a_LBL2_n_23 : std_logic;
  signal L1_L6a_LBL2_n_24, L1_L6a_LBL2_n_32, L1_L6a_c_rst_int, L1_L6a_eighty, L1_L6a_forty : std_logic;
  signal L1_L6a_hundredandtwenty, L1_L6a_sixty, L1_L6b_n_2, L1_L6b_n_3, L1_L6b_n_4 : std_logic;
  signal L1_L6b_n_5, L1_coin_present, L1_ghost1_ready, L1_ghost1_start, L1_ghost2_map_select : std_logic;
  signal L1_ghost2_start, L1_n_0, L1_n_1, L1_n_2, L1_n_3 : std_logic;
  signal L1_n_4, L1_n_5, L1_n_6, L1_n_7, L1_n_8 : std_logic;
  signal L1_n_9, L1_n_10, L1_n_11, L1_n_12, L1_n_13 : std_logic;
  signal L1_n_15, L1_n_16, L1_n_17, L1_n_18, L1_n_19 : std_logic;
  signal L1_n_20, L1_n_21, L1_n_22, L1_n_23, L1_n_24 : std_logic;
  signal L1_n_25, L1_n_26, L1_n_27, L1_n_28, L1_n_29 : std_logic;
  signal L1_n_30, L1_n_31, L1_n_32, L1_n_33, L1_n_34 : std_logic;
  signal L1_n_35, L1_n_36, L1_n_37, L1_n_38, L1_n_39 : std_logic;
  signal L1_n_40, L1_n_41, L1_n_42, L1_n_43, L1_n_44 : std_logic;
  signal L1_n_45, L1_n_46, L1_n_47, L1_n_48, L1_n_49 : std_logic;
  signal L1_n_50, L1_n_51, L1_n_52, L1_n_53, L1_n_54 : std_logic;
  signal L1_n_55, L1_n_56, L1_n_57, L1_n_58, L1_n_59 : std_logic;
  signal L1_n_60, L1_n_61, L1_n_62, L1_n_63, L1_n_64 : std_logic;
  signal L1_n_65, L1_n_66, L1_n_67, L1_n_68, L1_n_69 : std_logic;
  signal L1_n_70, L1_n_71, L1_n_72, L1_n_73, L1_n_74 : std_logic;
  signal L1_n_75, L1_n_76, L1_n_77, L1_n_78, L1_n_79 : std_logic;
  signal L1_n_80, L1_n_81, L1_n_82, L1_n_83, L1_n_84 : std_logic;
  signal L1_n_85, L1_n_86, L1_n_87, L1_n_88, L1_n_89 : std_logic;
  signal L1_n_90, L1_n_91, L1_n_92, L1_n_93, L1_n_94 : std_logic;
  signal L1_n_95, L1_n_96, L1_n_97, L1_n_98, L1_n_99 : std_logic;
  signal L1_n_100, L1_n_101, L1_n_102, L1_n_103, L1_n_104 : std_logic;
  signal L1_n_105, L1_n_106, L1_n_107, L1_n_108, L1_n_109 : std_logic;
  signal L1_n_110, L1_n_111, L1_n_112, L1_n_113, L1_n_114 : std_logic;
  signal L1_n_115, L1_n_116, L1_n_117, L1_n_118, L1_n_119 : std_logic;
  signal L1_n_120, L1_n_121, L1_n_122, L1_n_123, L1_n_124 : std_logic;
  signal L1_n_125, L1_n_126, L1_n_127, L1_n_128, L1_n_129 : std_logic;
  signal L1_n_130, L1_n_131, L1_n_132, L1_n_133, L1_n_134 : std_logic;
  signal L1_n_135, L1_n_136, L1_n_137, L1_n_138, L1_n_139 : std_logic;
  signal L1_n_140, L1_n_141, L1_n_142, L1_n_143, L1_n_144 : std_logic;
  signal L1_n_145, L1_n_146, L1_n_147, L1_n_148, L1_n_149 : std_logic;
  signal L1_n_150, L1_n_151, L1_n_152, L1_n_153, L1_n_154 : std_logic;
  signal L1_n_155, L1_n_156, L1_n_157, L1_n_158, L1_n_159 : std_logic;
  signal L1_n_160, L1_n_161, L1_n_162, L1_n_163, L1_n_164 : std_logic;
  signal L1_n_165, L1_n_166, L1_n_167, L1_n_168, L1_n_169 : std_logic;
  signal L1_n_170, L1_n_171, L1_n_172, L1_n_173, L1_n_174 : std_logic;
  signal L1_n_175, L1_n_176, L1_n_177, L1_n_178, L1_n_181 : std_logic;
  signal L1_n_182, L1_n_183, L1_n_184, L1_n_185, L1_n_186 : std_logic;
  signal L1_n_187, L1_n_188, L1_n_189, L1_n_190, L1_pacman_dead : std_logic;
  signal L1_pacman_map_select, L1_pacman_ready, L1_pacman_start, L1_pos_is_wall, L1_vc_pulse : std_logic;
  signal L1_write_coin, L1_zero_coins, L2_calc_start_internal, L2_dual_pixel_y, L2_en_county_go : std_logic;
  signal L2_en_county_score, L2_en_county_video, L2_en_current_block_horizontal_go, L2_en_current_block_horizontal_score, L2_en_current_block_horizontal_video : std_logic;
  signal L2_en_current_block_vertical, L2_en_dual_pixel_y_go, L2_en_dual_pixel_y_score, L2_en_dual_pixel_y_video, L2_gameovercontrol_n_2 : std_logic;
  signal L2_gameovercontrol_n_3, L2_gameovercontrol_n_4, L2_gameovercontrol_n_5, L2_gameovercontrol_n_6, L2_gameovercontrol_n_7 : std_logic;
  signal L2_gameovercontrol_n_8, L2_gameovercontrol_n_9, L2_gameovercontrol_n_10, L2_gameovercontrol_n_11, L2_gameovercontrol_n_12 : std_logic;
  signal L2_gameovercontrol_n_13, L2_gameovercontrol_n_14, L2_gameovercontrol_n_15, L2_gameovercontrol_n_16, L2_gameovercontrol_n_17 : std_logic;
  signal L2_gameovercontrol_n_18, L2_gameovercontrol_n_19, L2_gameovercontrol_n_20, L2_gameovercontrol_n_21, L2_gameovercontrol_n_22 : std_logic;
  signal L2_gameovercontrol_n_23, L2_gameovercontrol_n_24, L2_gameovercontrol_n_25, L2_gameovercontrol_n_26, L2_gameovercontrol_n_27 : std_logic;
  signal L2_gameovercontrol_n_28, L2_gameovercontrol_n_29, L2_gameovercontrol_n_30, L2_gameovercontrol_n_31, L2_gameovercontrol_n_32 : std_logic;
  signal L2_gameovercontrol_n_34, L2_gameovercontrol_n_35, L2_gameovercontrol_n_36, L2_gameovercontrol_n_37, L2_gameovercontrol_n_40 : std_logic;
  signal L2_gameovercontrol_n_41, L2_gameovercontrol_n_42, L2_gameovercontrol_n_43, L2_gameovercontrol_n_45, L2_gameovercontrol_n_46 : std_logic;
  signal L2_gameovercontrol_n_47, L2_gameovercontrol_n_48, L2_gameovercontrol_n_49, L2_gameovercontrol_n_50, L2_gameovercontrol_n_51 : std_logic;
  signal L2_gameovercontrol_n_52, L2_gameovercontrol_n_53, L2_gameovercontrol_n_54, L2_gameovercontrol_n_55, L2_gameovercontrol_n_56 : std_logic;
  signal L2_gameovercontrol_n_57, L2_gameovercontrol_n_58, L2_gameovercontrol_n_59, L2_gameovercontrol_n_60, L2_gameovercontrol_n_61 : std_logic;
  signal L2_gameovercontrol_n_62, L2_gameovercontrol_n_63, L2_gameovercontrol_n_64, L2_gameovercontrol_n_65, L2_gameovercontrol_n_66 : std_logic;
  signal L2_gameovercontrol_n_67, L2_gameovercontrol_n_68, L2_gameovercontrol_n_69, L2_gameovercontrol_n_70, L2_gameovercontrol_n_71 : std_logic;
  signal L2_gameovercontrol_n_72, L2_gameovercontrol_n_73, L2_gameovercontrol_n_74, L2_gameovercontrol_n_75, L2_gameovercontrol_n_76 : std_logic;
  signal L2_gameovercontrol_n_77, L2_gameovercontrol_n_78, L2_gameovercontrol_n_79, L2_gameovercontrol_n_80, L2_gameovercontrol_n_81 : std_logic;
  signal L2_gameovercontrol_n_82, L2_gameovercontrol_n_83, L2_gameovercontrol_n_84, L2_gameovercontrol_n_85, L2_gameovercontrol_n_86 : std_logic;
  signal L2_gameovercontrol_n_87, L2_gameovercontrol_n_88, L2_gameovercontrol_n_89, L2_gameovercontrol_n_90, L2_gameovercontrol_n_91 : std_logic;
  signal L2_gameovercontrol_n_92, L2_gameovercontrol_n_93, L2_gameovercontrol_n_94, L2_gameovercontrol_n_95, L2_gameovercontrol_n_96 : std_logic;
  signal L2_gameovercontrol_n_97, L2_gameovercontrol_n_98, L2_gameovercontrol_n_99, L2_gameovercontrol_n_100, L2_gameovercontrol_n_101 : std_logic;
  signal L2_gameovercontrol_n_102, L2_gameovercontrol_n_103, L2_gameovercontrol_n_104, L2_gameovercontrol_n_105, L2_gameovercontrol_n_106 : std_logic;
  signal L2_gameovercontrol_n_107, L2_gameovercontrol_n_108, L2_gameovercontrol_n_109, L2_gameovercontrol_n_110, L2_gameovercontrol_n_111 : std_logic;
  signal L2_gameovercontrol_n_112, L2_gameovercontrol_n_113, L2_gameovercontrol_n_114, L2_gameovercontrol_n_115, L2_gameovercontrol_n_116 : std_logic;
  signal L2_gameovercontrol_n_117, L2_gameovercontrol_n_118, L2_gameovercontrol_n_119, L2_gameovercontrol_n_120, L2_gameovercontrol_n_121 : std_logic;
  signal L2_gameovercontrol_n_122, L2_gameovercontrol_n_123, L2_gameovercontrol_n_124, L2_gameovercontrol_n_125, L2_gameovercontrol_n_126 : std_logic;
  signal L2_gameovercontrol_n_127, L2_gameovercontrol_n_128, L2_gameovercontrol_n_129, L2_gameovercontrol_n_131, L2_gameovercontrol_n_162 : std_logic;
  signal L2_gameovercontrol_n_163, L2_gameovercontrol_n_164, L2_gameovercontrol_n_165, L2_gameovercontrol_n_166, L2_gameovercontrol_n_976_BAR : std_logic;
  signal L2_gameovercontrol_row, L2_in_st_go_sel, L2_n_0, L2_n_1, L2_n_2 : std_logic;
  signal L2_n_3, L2_n_4, L2_n_5, L2_n_6, L2_n_7 : std_logic;
  signal L2_n_8, L2_n_9, L2_n_10, L2_n_11, L2_n_12 : std_logic;
  signal L2_n_13, L2_n_14, L2_n_15, L2_n_16, L2_n_17 : std_logic;
  signal L2_n_18, L2_n_19, L2_n_20, L2_n_21, L2_n_22 : std_logic;
  signal L2_n_23, L2_n_24, L2_n_25, L2_n_26, L2_n_27 : std_logic;
  signal L2_n_28, L2_n_29, L2_n_30, L2_n_31, L2_n_32 : std_logic;
  signal L2_n_33, L2_n_34, L2_n_35, L2_n_36, L2_n_37 : std_logic;
  signal L2_n_38, L2_n_39, L2_n_40, L2_n_41, L2_n_42 : std_logic;
  signal L2_n_43, L2_n_44, L2_n_45, L2_n_46, L2_n_47 : std_logic;
  signal L2_n_48, L2_n_49, L2_n_50, L2_n_51, L2_n_52 : std_logic;
  signal L2_n_53, L2_n_54, L2_n_55, L2_n_56, L2_n_57 : std_logic;
  signal L2_n_58, L2_n_59, L2_n_60, L2_n_61, L2_n_62 : std_logic;
  signal L2_n_63, L2_n_64, L2_n_65, L2_n_66, L2_n_67 : std_logic;
  signal L2_n_68, L2_n_69, L2_n_70, L2_n_71, L2_n_72 : std_logic;
  signal L2_n_73, L2_n_74, L2_n_75, L2_n_76, L2_n_77 : std_logic;
  signal L2_n_78, L2_n_79, L2_n_80, L2_n_81, L2_n_82 : std_logic;
  signal L2_n_83, L2_n_84, L2_n_85, L2_n_86, L2_n_87 : std_logic;
  signal L2_n_88, L2_n_89, L2_n_90, L2_n_91, L2_n_92 : std_logic;
  signal L2_n_93, L2_n_94, L2_n_95, L2_n_96, L2_n_97 : std_logic;
  signal L2_n_98, L2_n_99, L2_n_100, L2_n_101, L2_n_102 : std_logic;
  signal L2_n_103, L2_n_104, L2_n_105, L2_n_106, L2_n_107 : std_logic;
  signal L2_n_108, L2_n_109, L2_n_110, L2_n_111, L2_n_112 : std_logic;
  signal L2_n_113, L2_n_114, L2_n_115, L2_n_116, L2_n_117 : std_logic;
  signal L2_n_118, L2_n_119, L2_n_120, L2_n_121, L2_n_122 : std_logic;
  signal L2_n_123, L2_n_124, L2_n_125, L2_n_126, L2_n_127 : std_logic;
  signal L2_n_128, L2_n_129, L2_n_130, L2_n_131, L2_n_132 : std_logic;
  signal L2_n_133, L2_n_134, L2_n_135, L2_n_136, L2_n_137 : std_logic;
  signal L2_n_138, L2_n_139, L2_n_140, L2_n_141, L2_n_142 : std_logic;
  signal L2_n_143, L2_n_144, L2_n_145, L2_n_146, L2_n_147 : std_logic;
  signal L2_n_148, L2_n_149, L2_n_150, L2_n_151, L2_n_152 : std_logic;
  signal L2_n_153, L2_n_154, L2_n_155, L2_n_156, L2_n_157 : std_logic;
  signal L2_n_158, L2_n_159, L2_n_160, L2_n_161, L2_n_162 : std_logic;
  signal L2_n_163, L2_n_164, L2_n_165, L2_n_166, L2_n_167 : std_logic;
  signal L2_n_168, L2_n_169, L2_n_170, L2_n_171, L2_n_172 : std_logic;
  signal L2_n_173, L2_n_174, L2_n_175, L2_n_176, L2_n_177 : std_logic;
  signal L2_n_178, L2_n_179, L2_n_180, L2_n_181, L2_n_182 : std_logic;
  signal L2_n_183, L2_n_184, L2_n_185, L2_n_186, L2_n_187 : std_logic;
  signal L2_n_188, L2_n_189, L2_n_190, L2_n_191, L2_n_192 : std_logic;
  signal L2_n_193, L2_n_194, L2_n_195, L2_n_196, L2_n_197 : std_logic;
  signal L2_n_198, L2_n_199, L2_n_200, L2_n_201, L2_n_202 : std_logic;
  signal L2_n_203, L2_n_204, L2_n_205, L2_n_206, L2_n_207 : std_logic;
  signal L2_n_208, L2_n_209, L2_n_210, L2_n_211, L2_n_212 : std_logic;
  signal L2_n_213, L2_n_214, L2_n_215, L2_n_216, L2_n_217 : std_logic;
  signal L2_n_218, L2_n_219, L2_n_220, L2_n_221, L2_n_222 : std_logic;
  signal L2_n_223, L2_n_224, L2_n_225, L2_n_226, L2_n_227 : std_logic;
  signal L2_n_228, L2_n_229, L2_n_230, L2_n_231, L2_n_232 : std_logic;
  signal L2_n_233, L2_n_234, L2_n_235, L2_n_236, L2_n_237 : std_logic;
  signal L2_n_238, L2_n_239, L2_n_240, L2_n_241, L2_n_242 : std_logic;
  signal L2_n_243, L2_n_244, L2_n_245, L2_n_246, L2_n_247 : std_logic;
  signal L2_n_248, L2_n_249, L2_n_250, L2_n_251, L2_n_252 : std_logic;
  signal L2_n_253, L2_n_254, L2_n_255, L2_n_256, L2_n_257 : std_logic;
  signal L2_n_258, L2_n_259, L2_n_260, L2_n_261, L2_n_262 : std_logic;
  signal L2_n_263, L2_n_264, L2_n_265, L2_n_266, L2_n_267 : std_logic;
  signal L2_n_268, L2_n_269, L2_n_270, L2_n_271, L2_n_272 : std_logic;
  signal L2_n_273, L2_n_274, L2_n_275, L2_n_276, L2_n_277 : std_logic;
  signal L2_n_278, L2_n_279, L2_n_280, L2_n_281, L2_n_282 : std_logic;
  signal L2_n_283, L2_n_284, L2_n_285, L2_n_286, L2_n_287 : std_logic;
  signal L2_n_288, L2_n_289, L2_n_290, L2_n_291, L2_n_292 : std_logic;
  signal L2_n_293, L2_n_294, L2_n_295, L2_n_296, L2_n_297 : std_logic;
  signal L2_n_298, L2_n_299, L2_n_300, L2_n_301, L2_n_302 : std_logic;
  signal L2_n_303, L2_n_304, L2_n_305, L2_n_306, L2_n_307 : std_logic;
  signal L2_n_308, L2_n_309, L2_n_310, L2_n_311, L2_n_312 : std_logic;
  signal L2_n_313, L2_n_314, L2_n_315, L2_n_316, L2_n_317 : std_logic;
  signal L2_n_318, L2_n_319, L2_n_320, L2_n_321, L2_n_322 : std_logic;
  signal L2_n_323, L2_n_324, L2_n_325, L2_n_326, L2_n_327 : std_logic;
  signal L2_n_328, L2_n_329, L2_n_330, L2_n_331, L2_n_332 : std_logic;
  signal L2_n_333, L2_n_334, L2_n_335, L2_n_336, L2_n_337 : std_logic;
  signal L2_n_338, L2_n_339, L2_n_340, L2_n_341, L2_n_342 : std_logic;
  signal L2_n_343, L2_n_344, L2_n_345, L2_n_346, L2_n_347 : std_logic;
  signal L2_n_348, L2_n_349, L2_n_350, L2_n_351, L2_n_352 : std_logic;
  signal L2_n_353, L2_n_354, L2_n_355, L2_n_356, L2_n_357 : std_logic;
  signal L2_n_358, L2_n_359, L2_n_360, L2_n_361, L2_n_362 : std_logic;
  signal L2_n_363, L2_n_364, L2_n_365, L2_n_366, L2_n_367 : std_logic;
  signal L2_n_368, L2_n_369, L2_n_370, L2_n_371, L2_n_372 : std_logic;
  signal L2_n_373, L2_n_374, L2_n_375, L2_n_376, L2_n_377 : std_logic;
  signal L2_n_378, L2_n_379, L2_n_380, L2_n_381, L2_n_382 : std_logic;
  signal L2_n_383, L2_n_384, L2_n_385, L2_n_386, L2_n_387 : std_logic;
  signal L2_n_388, L2_n_389, L2_n_390, L2_n_391, L2_n_392 : std_logic;
  signal L2_n_393, L2_n_394, L2_n_395, L2_n_396, L2_n_397 : std_logic;
  signal L2_n_398, L2_n_399, L2_n_400, L2_n_401, L2_n_402 : std_logic;
  signal L2_n_403, L2_n_404, L2_n_405, L2_n_406, L2_n_407 : std_logic;
  signal L2_n_408, L2_n_409, L2_n_410, L2_n_411, L2_n_412 : std_logic;
  signal L2_n_413, L2_n_414, L2_n_415, L2_n_416, L2_n_417 : std_logic;
  signal L2_n_418, L2_n_419, L2_n_420, L2_n_421, L2_n_422 : std_logic;
  signal L2_n_423, L2_n_424, L2_n_425, L2_n_426, L2_n_427 : std_logic;
  signal L2_n_428, L2_n_429, L2_n_430, L2_n_431, L2_n_432 : std_logic;
  signal L2_n_433, L2_n_434, L2_n_435, L2_n_436, L2_n_437 : std_logic;
  signal L2_n_438, L2_n_439, L2_n_440, L2_n_441, L2_n_442 : std_logic;
  signal L2_n_443, L2_n_444, L2_n_445, L2_n_446, L2_n_447 : std_logic;
  signal L2_n_448, L2_n_449, L2_n_450, L2_n_451, L2_n_452 : std_logic;
  signal L2_n_453, L2_n_454, L2_n_455, L2_n_456, L2_n_457 : std_logic;
  signal L2_n_458, L2_n_459, L2_n_460, L2_n_461, L2_n_462 : std_logic;
  signal L2_n_463, L2_n_464, L2_n_465, L2_n_466, L2_n_467 : std_logic;
  signal L2_n_468, L2_n_469, L2_n_470, L2_n_471, L2_n_472 : std_logic;
  signal L2_n_473, L2_n_474, L2_n_475, L2_n_476, L2_n_477 : std_logic;
  signal L2_n_478, L2_n_479, L2_n_480, L2_n_481, L2_n_482 : std_logic;
  signal L2_n_483, L2_n_484, L2_n_485, L2_n_486, L2_n_487 : std_logic;
  signal L2_n_488, L2_n_489, L2_n_490, L2_n_491, L2_n_492 : std_logic;
  signal L2_n_493, L2_n_494, L2_n_495, L2_n_496, L2_n_497 : std_logic;
  signal L2_n_498, L2_n_499, L2_n_500, L2_n_501, L2_n_502 : std_logic;
  signal L2_n_503, L2_n_504, L2_n_505, L2_n_506, L2_n_507 : std_logic;
  signal L2_n_508, L2_n_509, L2_n_510, L2_n_511, L2_n_512 : std_logic;
  signal L2_n_513, L2_n_514, L2_n_515, L2_n_516, L2_n_517 : std_logic;
  signal L2_n_518, L2_n_519, L2_n_521, L2_n_522, L2_n_523 : std_logic;
  signal L2_n_524, L2_n_525, L2_n_526, L2_n_527, L2_n_528 : std_logic;
  signal L2_n_529, L2_n_530, L2_n_531, L2_n_532, L2_n_533 : std_logic;
  signal L2_n_534, L2_n_535, L2_n_536, L2_n_537, L2_n_538 : std_logic;
  signal L2_n_539, L2_n_540, L2_n_541, L2_n_542, L2_n_543 : std_logic;
  signal L2_n_544, L2_n_545, L2_n_546, L2_n_547, L2_n_548 : std_logic;
  signal L2_n_549, L2_n_550, L2_n_551, L2_n_552, L2_reset_county_go : std_logic;
  signal L2_reset_county_score, L2_reset_county_video, L2_reset_current_block_horizontal_go, L2_reset_current_block_horizontal_score, L2_reset_current_block_horizontal_video : std_logic;
  signal L2_reset_current_block_vertical, L2_reset_dual_pixel_y_go, L2_reset_dual_pixel_y_score, L2_reset_dual_pixel_y_video, L2_score_L2_n_0 : std_logic;
  signal L2_score_L2_n_1, L2_score_L2_n_4, L2_score_L2_n_5, L2_score_L2_n_6, L2_score_L2_n_7 : std_logic;
  signal L2_score_L2_n_8, L2_score_L2_n_9, L2_score_L2_n_10, L2_score_L2_n_11, L2_score_L2_n_12 : std_logic;
  signal L2_score_L2_n_13, L2_score_L2_n_14, L2_score_L2_n_15, L2_score_L2_n_16, L2_score_L2_n_17 : std_logic;
  signal L2_score_L2_n_18, L2_score_L2_n_19, L2_score_L2_n_20, L2_score_L2_n_21, L2_score_L2_n_22 : std_logic;
  signal L2_score_L2_n_23, L2_score_L2_n_24, L2_score_L2_n_25, L2_score_L2_n_26, L2_score_L2_n_27 : std_logic;
  signal L2_score_L2_n_28, L2_score_L2_n_29, L2_score_L2_n_30, L2_score_L2_n_31, L2_score_L2_n_32 : std_logic;
  signal L2_score_L2_n_33, L2_score_L2_n_34, L2_score_L2_n_35, L2_score_L2_n_36, L2_score_L2_n_37 : std_logic;
  signal L2_score_L2_n_38, L2_score_L2_n_39, L2_score_L2_n_40, L2_score_L2_n_41, L2_score_L2_n_42 : std_logic;
  signal L2_score_L2_n_43, L2_score_L2_n_44, L2_score_L2_n_45, L2_score_L2_n_46, L2_score_L2_n_47 : std_logic;
  signal L2_score_L2_n_48, L2_score_L2_n_49, L2_score_L2_n_50, L2_score_L2_n_51, L2_score_L2_n_52 : std_logic;
  signal L2_score_L2_n_53, L2_score_L2_n_54, L2_score_L2_n_55, L2_score_L2_n_56, L2_score_L2_n_57 : std_logic;
  signal L2_score_L2_n_58, L2_score_L3_n_0, L2_score_L3_n_1, L2_score_L3_n_2, L2_score_L3_n_3 : std_logic;
  signal L2_score_L3_n_4, L2_score_L3_n_5, L2_score_L3_n_6, L2_score_L3_n_7, L2_score_L3_n_8 : std_logic;
  signal L2_score_L3_n_9, L2_score_L3_n_10, L2_score_L3_n_12, L2_score_L3_n_13, L2_score_L3_n_14 : std_logic;
  signal L2_score_L3_n_15, L2_score_L3_n_16, L2_score_L3_n_17, L2_score_L3_n_18, L2_score_L3_n_19 : std_logic;
  signal L2_score_L3_n_20, L2_score_L3_n_21, L2_score_L3_n_22, L2_score_L3_n_23, L2_score_L3_n_24 : std_logic;
  signal L2_score_L3_n_25, L2_score_L3_n_26, L2_score_L3_n_27, L2_score_L3_n_28, L2_score_L3_n_29 : std_logic;
  signal L2_score_L3_n_30, L2_score_L3_n_31, L2_score_L3_n_32, L2_score_L3_n_33, L2_score_L3_n_34 : std_logic;
  signal L2_score_L3_n_35, L2_score_L3_n_36, L2_score_L3_n_37, L2_score_L3_n_38, L2_score_L3_n_39 : std_logic;
  signal L2_score_L3_n_40, L2_score_L3_n_41, L2_score_L3_n_42, L2_score_L3_n_43, L2_score_L3_n_44 : std_logic;
  signal L2_score_L3_n_45, L2_score_L3_n_46, L2_score_L3_n_47, L2_score_L3_n_48, L2_score_L3_n_49 : std_logic;
  signal L2_score_L3_n_50, L2_score_L3_n_51, L2_score_L3_n_52, L2_score_L3_n_53, L2_score_L3_n_54 : std_logic;
  signal L2_score_L3_n_55, L2_score_L3_n_56, L2_score_L3_n_57, L2_score_L3_n_58, L2_score_L3_n_59 : std_logic;
  signal L2_score_L3_n_60, L2_score_L3_n_61, L2_score_L3_n_62, L2_score_L3_n_63, L2_score_L3_n_64 : std_logic;
  signal L2_score_L3_n_65, L2_score_L3_n_66, L2_score_L3_n_67, L2_score_L3_n_68, L2_score_L3_n_69 : std_logic;
  signal L2_score_L3_n_70, L2_score_L3_n_71, L2_score_L3_n_72, L2_score_L3_n_73, L2_score_L3_n_74 : std_logic;
  signal L2_score_L3_n_75, L2_score_L3_n_76, L2_score_L3_n_77, L2_score_L3_n_78, L2_score_L3_n_79 : std_logic;
  signal L2_score_L3_n_80, L2_score_L3_n_81, L2_score_L3_n_83, L2_score_L3_n_84, L2_score_L3_n_87 : std_logic;
  signal L2_score_L3_n_88, L2_score_L3_n_89, L2_score_L3_n_90, L2_score_L3_n_91, L2_score_L3_n_93 : std_logic;
  signal L2_score_L3_n_94, L2_score_L3_n_95, L2_score_L3_n_135, L2_score_reset_or, L2_screencontrol_go : std_logic;
  signal L2_screencontrol_n_58, L2_screencontrol_n_66, L2_shift_L11_n_0, L2_shift_L11_n_1, L2_shift_L11_n_2 : std_logic;
  signal L2_shift_L11_n_3, L2_shift_L11_n_4, L2_shift_L11_n_5, L2_shift_L11_n_6, L2_shift_L11_n_7 : std_logic;
  signal L2_shift_L11_n_8, L2_shift_L11_n_9, L2_shift_L11_n_10, L2_shift_L11_n_11, L2_shift_L11_n_12 : std_logic;
  signal L2_shift_L11_n_13, L2_shift_L11_n_14, L2_shift_L11_n_15, L2_shift_L11_n_16, L2_shift_L11_n_17 : std_logic;
  signal L2_shift_L11_n_18, L2_shift_L11_n_19, L2_shift_L11_n_20, L2_shift_L11_n_21, L2_shift_L11_n_22 : std_logic;
  signal L2_shift_L11_n_23, L2_shift_L11_n_24, L2_shift_L11_n_25, L2_shift_L11_n_26, L2_shift_L11_n_27 : std_logic;
  signal L2_shift_L11_n_28, L2_shift_L11_n_29, L2_shift_L11_n_30, L2_shift_L11_n_31, L2_shift_L11_n_32 : std_logic;
  signal L2_shift_L11_n_33, L2_shift_L11_n_34, L2_shift_L11_n_35, L2_shift_L11_n_36, L2_shift_L11_n_37 : std_logic;
  signal L2_shift_L11_n_38, L2_shift_L11_n_39, L2_shift_L11_n_40, L2_shift_L11_n_41, L2_shift_L11_n_42 : std_logic;
  signal L2_shift_L11_n_43, L2_shift_L11_n_44, L2_shift_L11_n_45, L2_shift_L11_n_46, L2_shift_L11_n_47 : std_logic;
  signal L2_shift_L11_n_48, L2_shift_L11_n_49, L2_shift_L11_n_50, L2_shift_L11_n_51, L2_shift_L11_n_52 : std_logic;
  signal L2_shift_L11_n_53, L2_shift_L11_n_54, L2_shift_L11_n_55, L2_shift_L11_n_56, L2_shift_L11_n_57 : std_logic;
  signal L2_shift_L11_n_58, L2_shift_L11_n_59, L2_shift_L11_n_60, L2_shift_L11_n_61, L2_shift_L11_n_62 : std_logic;
  signal L2_shift_L11_n_63, L2_shift_L11_n_64, L2_shift_L11_n_65, L2_shift_L11_n_66, L2_shift_L11_n_67 : std_logic;
  signal L2_shift_L11_n_68, L2_shift_L11_n_69, L2_shift_L11_n_70, L2_shift_L11_n_71, L2_shift_L11_n_72 : std_logic;
  signal L2_shift_L11_n_73, L2_shift_L11_n_74, L2_shift_L11_n_75, L2_shift_L11_n_76, L2_shift_L11_n_77 : std_logic;
  signal L2_shift_L11_n_78, L2_shift_L11_n_79, L2_shift_L11_n_80, L2_shift_L11_n_81, L2_shift_L11_n_82 : std_logic;
  signal L2_shift_L11_n_83, L2_shift_L11_n_84, L2_shift_L11_n_85, L2_shift_L11_n_86, L2_shift_L11_n_87 : std_logic;
  signal L2_shift_L11_n_88, L2_shift_L11_n_89, L2_shift_L11_n_90, L2_shift_L11_n_91, L2_shift_L11_n_92 : std_logic;
  signal L2_shift_L11_n_93, L2_shift_L11_n_94, L2_shift_L11_n_95, L2_shift_L11_n_96, L2_shift_L11_n_97 : std_logic;
  signal L2_shift_L11_n_98, L2_shift_L11_n_99, L2_shift_L11_n_100, L2_shift_L11_n_101, L2_shift_L11_n_102 : std_logic;
  signal L2_shift_L11_n_103, L2_shift_L11_n_104, L2_shift_L11_n_105, L2_shift_L11_n_106, L2_shift_L11_n_107 : std_logic;
  signal L2_shift_L11_n_108, L2_shift_L11_n_109, L2_shift_L11_n_110, L2_shift_L11_n_111, L2_shift_L11_n_112 : std_logic;
  signal L2_shift_L11_n_113, L2_shift_L11_n_114, L2_shift_L11_n_115, L2_shift_L11_n_116, L2_shift_L11_n_118 : std_logic;
  signal L2_shift_L11_n_119, L2_shift_L11_n_120, L2_shift_L11_n_121, L2_shift_L11_n_122, L2_shift_L11_n_123 : std_logic;
  signal L2_shift_L11_n_124, L2_shift_L11_n_125, L2_shift_L11_n_126, L2_shift_L11_n_127, L2_shift_L11_n_128 : std_logic;
  signal L2_shift_L11_n_129, L2_shift_L11_n_130, L2_shift_L11_n_131, L2_shift_L11_n_132, L2_shift_L11_n_133 : std_logic;
  signal L2_shift_L11_n_134, L2_shift_L11_n_135, L2_shift_L11_n_136, L2_shift_L11_n_137, L2_shift_L11_n_138 : std_logic;
  signal L2_shift_L11_n_139, L2_shift_L11_n_140, L2_shift_L11_n_141, L2_shift_L11_n_142, L2_shift_L11_n_143 : std_logic;
  signal L2_shift_L11_n_144, L2_shift_L11_n_146, L2_shift_L11_n_147, L2_shift_L11_n_148, L2_shift_L11_n_149 : std_logic;
  signal L2_shift_L11_n_150, L2_shift_L11_n_151, L2_shift_L11_n_152, L2_shift_L11_n_153, L2_shift_L11_n_154 : std_logic;
  signal L2_shift_L11_n_155, L2_shift_L11_n_156, L2_shift_L11_n_157, L2_shift_L11_n_158, L2_shift_L11_n_159 : std_logic;
  signal L2_shift_L11_n_160, L2_shift_L11_n_161, L2_shift_L11_n_162, L2_shift_L11_n_163, L2_shift_L11_n_164 : std_logic;
  signal L2_shift_L11_n_165, L2_shift_L11_n_166, L2_shift_L11_n_167, L2_shift_L11_n_168, L2_shift_L11_n_169 : std_logic;
  signal L2_shift_L11_n_170, L2_shift_L11_n_171, L2_shift_L11_n_172, L2_shift_L11_n_173, L2_shift_L11_n_174 : std_logic;
  signal L2_shift_L11_n_175, L2_shift_L11_n_176, L2_shift_L11_n_177, L2_shift_L11_n_178, L2_shift_L11_n_179 : std_logic;
  signal L2_shift_L11_n_180, L2_shift_L11_n_181, L2_shift_L11_n_182, L2_shift_L11_n_183, L2_shift_L11_n_184 : std_logic;
  signal L2_shift_L11_n_185, L2_shift_L11_n_186, L2_shift_L11_n_187, L2_shift_L11_n_188, L2_shift_L11_n_189 : std_logic;
  signal L2_shift_L11_n_190, L2_shift_L11_n_191, L2_shift_L11_n_192, L2_shift_L11_n_193, L2_shift_L11_n_194 : std_logic;
  signal L2_shift_L11_n_195, L2_shift_L11_n_196, L2_shift_L11_n_197, L2_shift_L11_n_198, L2_shift_L11_n_199 : std_logic;
  signal L2_shift_L11_n_200, L2_shift_L11_n_201, L2_shift_L11_n_202, L2_shift_L11_n_203, L2_shift_L11_n_204 : std_logic;
  signal L2_shift_L11_n_205, L2_shift_L11_n_206, L2_shift_L11_n_207, L2_shift_L11_n_208, L2_shift_L11_n_209 : std_logic;
  signal L2_shift_L11_n_210, L2_shift_L11_n_211, L2_shift_L11_n_212, L2_shift_L11_n_213, L2_shift_L11_n_214 : std_logic;
  signal L2_shift_L11_n_215, L2_shift_L11_n_216, L2_shift_L11_n_217, L2_shift_L11_n_218, L2_shift_L11_n_219 : std_logic;
  signal L2_shift_L11_n_220, L2_shift_L11_n_221, L2_shift_L11_n_222, L2_shift_L11_n_223, L2_shift_L11_n_224 : std_logic;
  signal L2_shift_L11_n_225, L2_shift_L11_n_226, L2_shift_L11_n_227, L2_shift_L11_n_228, L2_shift_L11_n_229 : std_logic;
  signal L2_shift_L11_n_230, L2_shift_L11_n_231, L2_shift_L11_n_232, L2_shift_L11_n_233, L2_shift_L11_n_234 : std_logic;
  signal L2_shift_L11_n_235, L2_shift_L11_n_236, L2_shift_L11_n_237, L2_shift_L11_n_238, L2_shift_L11_n_239 : std_logic;
  signal L2_shift_L11_n_240, L2_shift_L11_n_241, L2_shift_L11_n_242, L2_shift_L11_n_243, L2_shift_L11_n_244 : std_logic;
  signal L2_shift_L11_n_245, L2_shift_L11_n_246, L2_shift_L11_n_247, L2_shift_L11_n_248, L2_shift_L11_n_249 : std_logic;
  signal L2_shift_L11_n_250, L2_shift_L11_n_251, L2_shift_L11_n_252, L2_shift_L11_n_253, L2_shift_L11_n_254 : std_logic;
  signal L2_shift_L11_n_255, L2_shift_L11_n_256, L2_shift_L11_n_257, L2_shift_L11_n_258, L2_shift_L11_n_259 : std_logic;
  signal L2_shift_L11_n_260, L2_shift_L11_n_261, L2_shift_L11_n_262, L2_shift_L11_n_263, L2_shift_L11_n_264 : std_logic;
  signal L2_shift_L11_n_265, L2_shift_L11_n_266, L2_shift_L11_n_267, L2_shift_L11_n_268, L2_shift_L11_n_269 : std_logic;
  signal L2_shift_L11_n_270, L2_shift_L11_n_271, L2_shift_L11_n_272, L2_shift_L11_n_273, L2_shift_L11_n_274 : std_logic;
  signal L2_shift_L11_n_275, L2_shift_L11_n_276, L2_shift_L11_n_277, L2_shift_L11_n_278, L2_shift_L11_n_279 : std_logic;
  signal L2_shift_L11_n_280, L2_shift_L11_n_281, L2_shift_L11_n_282, L2_shift_L11_n_283, L2_shift_L11_n_284 : std_logic;
  signal L2_shift_L11_n_285, L2_shift_L11_n_286, L2_shift_L11_n_287, L2_shift_L11_n_288, L2_shift_L11_n_289 : std_logic;
  signal L2_shift_L11_n_290, L2_shift_L11_n_292, L2_shift_L11_n_293, L2_shift_L11_n_294, L2_shift_L11_n_295 : std_logic;
  signal L2_shift_L11_n_296, L2_shift_L11_n_297, L2_shift_L11_n_298, L2_shift_L11_n_299, L2_shift_L11_n_302 : std_logic;
  signal L2_shift_L11_n_303, L2_shift_L11_n_304, L2_shift_L11_n_305, L2_shift_L11_n_306, L2_shift_L11_n_307 : std_logic;
  signal L2_shift_L11_n_308, L2_shift_L11_n_309, L2_shift_L11_n_310, L2_shift_L11_n_311, L2_shift_L11_n_312 : std_logic;
  signal L2_shift_L11_n_313, L2_shift_L11_n_314, L2_shift_L11_n_315, L2_shift_L11_n_316, L2_shift_L11_n_317 : std_logic;
  signal L2_shift_L11_n_318, L2_shift_L11_n_319, L2_shift_L11_n_320, L2_shift_L11_n_321, L2_shift_L11_n_322 : std_logic;
  signal L2_shift_L11_n_323, L2_shift_L11_n_324, L2_shift_L11_n_325, L2_shift_L11_n_326, L2_shift_L11_n_327 : std_logic;
  signal L2_shift_L11_n_328, L2_shift_L11_n_329, L2_shift_L11_n_330, L2_shift_L11_n_331, L2_shift_L11_n_332 : std_logic;
  signal L2_shift_L11_n_333, L2_shift_L11_n_334, L2_shift_L11_n_335, L2_shift_L11_n_336, L2_shift_L11_n_337 : std_logic;
  signal L2_shift_L11_n_399, L2_shift_L11_n_403, L2_shift_L11_n_405, L2_shift_L11_n_406, L2_shift_L11_n_407 : std_logic;
  signal L2_shift_L21_n_0, L2_shift_L21_n_1, L2_shift_L21_n_2, L2_shift_L21_n_3, L2_shift_L21_n_4 : std_logic;
  signal L2_shift_L21_n_5, L2_shift_L21_n_6, L2_shift_L21_n_7, L2_shift_L21_n_8, L2_shift_L21_n_9 : std_logic;
  signal L2_shift_L21_n_10, L2_shift_L23_n_1, L2_shift_L23_n_2, L2_shift_L23_n_3, L2_shift_L23_n_4 : std_logic;
  signal L2_shift_L23_n_5, L2_shift_L23_n_6, L2_shift_L23_n_7, L2_shift_L23_n_8, L2_shift_L23_n_9 : std_logic;
  signal L2_shift_L23_n_10, L2_shift_L23_n_11, L2_shift_L23_n_12, L2_shift_L23_n_13, L2_shift_L23_n_14 : std_logic;
  signal L2_shift_L23_n_15, L2_shift_L23_n_16, L2_shift_L23_n_17, L2_shift_L23_n_18, L2_shift_L23_n_19 : std_logic;
  signal L2_shift_L23_n_20, L2_shift_L23_n_21, L2_shift_L23_n_22, L2_shift_L23_n_23, L2_shift_L23_n_24 : std_logic;
  signal L2_shift_L23_n_25, L2_shift_L23_n_26, L2_shift_L23_n_27, L2_shift_L23_n_28, L2_shift_L23_n_29 : std_logic;
  signal L2_shift_L23_n_30, L2_shift_L23_n_31, L2_shift_L23_n_32, L2_shift_L23_n_33, L2_shift_L23_n_34 : std_logic;
  signal L2_shift_L23_n_35, L2_shift_L23_n_36, L2_shift_L23_n_37, L2_shift_L23_n_38, L2_shift_L23_n_39 : std_logic;
  signal L2_shift_L23_n_40, L2_shift_L23_n_41, L2_shift_L23_n_42, L2_shift_L23_n_43, L2_shift_L23_n_44 : std_logic;
  signal L2_shift_L23_n_45, L2_shift_L23_n_46, L2_shift_L23_n_47, L2_shift_L23_n_48, L2_shift_L23_n_49 : std_logic;
  signal L2_shift_L23_n_50, L2_shift_L23_n_51, L2_shift_L23_n_52, L2_shift_L23_n_53, L2_shift_L23_n_54 : std_logic;
  signal L2_shift_L23_n_55, L2_shift_L23_n_56, L2_shift_L23_n_57, L2_shift_L23_n_58, L2_shift_L23_n_59 : std_logic;
  signal L2_shift_L23_n_60, L2_shift_L23_n_61, L2_shift_L23_n_62, L2_shift_L23_n_63, L2_shift_L23_n_64 : std_logic;
  signal L2_shift_L23_n_65, L2_shift_L23_n_66, L2_shift_L23_n_67, L2_shift_L23_n_68, L2_shift_L23_n_69 : std_logic;
  signal L2_shift_L23_n_70, L2_shift_L23_n_71, L2_shift_L23_n_72, L2_shift_L23_n_73, L2_shift_L23_n_74 : std_logic;
  signal L2_shift_L23_n_75, L2_shift_L23_n_76, L2_shift_L23_n_77, L2_shift_L23_n_78, L2_shift_L23_n_79 : std_logic;
  signal L2_shift_L23_n_80, L2_shift_L23_n_81, L2_shift_L23_n_82, L2_shift_L23_n_83, L2_shift_L23_n_84 : std_logic;
  signal L2_shift_L23_n_85, L2_shift_L23_n_86, L2_shift_L23_n_87, L2_shift_L23_n_88, L2_shift_L23_n_89 : std_logic;
  signal L2_shift_L23_n_90, L2_shift_L23_n_91, L2_shift_L23_n_92, L2_shift_L23_n_93, L2_shift_L23_n_94 : std_logic;
  signal L2_shift_L23_n_95, L2_shift_L23_n_96, L2_shift_L23_n_97, L2_shift_L23_n_98, L2_shift_L23_n_99 : std_logic;
  signal L2_shift_L23_n_100, L2_shift_L23_n_101, L2_shift_L23_n_102, L2_shift_L23_n_103, L2_shift_L23_n_104 : std_logic;
  signal L2_shift_L23_n_105, L2_shift_L23_n_106, L2_shift_L23_n_107, L2_shift_L23_n_108, L2_shift_L23_n_109 : std_logic;
  signal L2_shift_L23_n_110, L2_shift_L23_n_111, L2_shift_L23_n_112, L2_shift_L23_n_113, L2_shift_L23_n_114 : std_logic;
  signal L2_shift_L23_n_115, L2_shift_L23_n_116, L2_shift_L23_n_117, L2_shift_L23_n_118, L2_shift_L23_n_119 : std_logic;
  signal L2_shift_L23_n_120, L2_shift_L23_n_121, L2_shift_L23_n_122, L2_shift_L23_n_123, L2_shift_L23_n_124 : std_logic;
  signal L2_shift_L23_n_125, L2_shift_L23_n_126, L2_shift_L23_n_127, L2_shift_L23_n_128, L2_shift_L23_n_129 : std_logic;
  signal L2_shift_L23_n_131, L2_shift_L23_n_132, L2_shift_L23_n_133, L2_shift_L23_n_134, L2_shift_L23_n_135 : std_logic;
  signal L2_shift_L23_n_136, L2_shift_L23_n_137, L2_shift_L23_n_138, L2_shift_L23_n_139, L2_shift_L23_n_140 : std_logic;
  signal L2_shift_L23_n_141, L2_shift_L23_n_142, L2_shift_L23_n_143, L2_shift_L23_n_144, L2_shift_L23_n_145 : std_logic;
  signal L2_shift_L23_n_146, L2_shift_L23_n_148, L2_shift_L23_n_149, L2_shift_L23_n_150, L2_shift_L23_n_151 : std_logic;
  signal L2_shift_L23_n_152, L2_shift_L23_n_154, L2_shift_L23_n_155, L2_shift_L23_n_156, L2_shift_L23_n_157 : std_logic;
  signal L2_shift_L23_n_158, L2_shift_L23_n_159, L2_shift_L23_n_160, L2_shift_L23_n_161, L2_shift_L23_n_162 : std_logic;
  signal L2_shift_L23_n_163, L2_shift_L23_n_164, L2_shift_L23_n_165, L2_shift_L23_n_166, L2_shift_L23_n_167 : std_logic;
  signal L2_shift_L23_n_168, L2_shift_L23_n_169, L2_shift_L23_n_170, L2_shift_L23_n_171, L2_shift_L23_n_172 : std_logic;
  signal L2_shift_L23_n_173, L2_shift_L23_n_174, L2_shift_L23_n_175, L2_shift_L23_n_176, L2_shift_L23_n_177 : std_logic;
  signal L2_shift_L23_n_178, L2_shift_L23_n_179, L2_shift_L23_n_180, L2_shift_L23_n_181, L2_shift_L23_n_182 : std_logic;
  signal L2_shift_L23_n_183, L2_shift_L23_n_184, L2_shift_L23_n_185, L2_shift_L23_n_186, L2_shift_L23_n_187 : std_logic;
  signal L2_shift_L23_n_188, L2_shift_L23_n_189, L2_shift_L23_n_190, L2_shift_L23_n_191, L2_shift_L23_n_192 : std_logic;
  signal L2_shift_L23_n_193, L2_shift_L23_n_194, L2_shift_L23_n_195, L2_shift_L23_n_196, L2_shift_L23_n_197 : std_logic;
  signal L2_shift_L23_n_198, L2_shift_L23_n_199, L2_shift_L23_n_200, L2_shift_L23_n_201, L2_shift_L23_n_202 : std_logic;
  signal L2_shift_L23_n_203, L2_shift_L23_n_204, L2_shift_L23_n_205, L2_shift_L23_n_206, L2_shift_L23_n_207 : std_logic;
  signal L2_shift_L23_n_208, L2_shift_L23_n_209, L2_shift_L23_n_210, L2_shift_L23_n_211, L2_shift_L23_n_212 : std_logic;
  signal L2_shift_L23_n_213, L2_shift_L23_n_214, L2_shift_L23_n_215, L2_shift_L23_n_216, L2_shift_L23_n_217 : std_logic;
  signal L2_shift_L23_n_218, L2_shift_L23_n_219, L2_shift_L23_n_220, L2_shift_L23_n_221, L2_shift_L23_n_222 : std_logic;
  signal L2_shift_L23_n_223, L2_shift_L23_n_224, L2_shift_L23_n_225, L2_shift_L23_n_226, L2_shift_L23_n_227 : std_logic;
  signal L2_shift_L23_n_228, L2_shift_L23_n_229, L2_shift_L23_n_230, L2_shift_L23_n_231, L2_shift_L23_n_232 : std_logic;
  signal L2_shift_L23_n_233, L2_shift_L23_n_234, L2_shift_L23_n_235, L2_shift_L23_n_236, L2_shift_L23_n_237 : std_logic;
  signal L2_shift_L23_n_238, L2_shift_L23_n_239, L2_shift_L23_n_240, L2_shift_L23_n_241, L2_shift_L23_n_242 : std_logic;
  signal L2_shift_L23_n_243, L2_shift_L23_n_244, L2_shift_L23_n_245, L2_shift_L23_n_246, L2_shift_L23_n_247 : std_logic;
  signal L2_shift_L23_n_248, L2_shift_L23_n_249, L2_shift_L23_n_250, L2_shift_L23_n_251, L2_shift_L23_n_252 : std_logic;
  signal L2_shift_L23_n_253, L2_shift_L23_n_254, L2_shift_L23_n_255, L2_shift_L23_n_256, L2_shift_L23_n_257 : std_logic;
  signal L2_shift_L23_n_258, L2_shift_L23_n_259, L2_shift_L23_n_260, L2_shift_L23_n_261, L2_shift_L23_n_262 : std_logic;
  signal L2_shift_L23_n_263, L2_shift_L23_n_264, L2_shift_L23_n_265, L2_shift_L23_n_267, L2_shift_L23_n_268 : std_logic;
  signal L2_shift_L23_n_269, L2_shift_L23_n_271, L2_shift_L23_n_272, L2_shift_L23_n_273, L2_shift_L23_n_274 : std_logic;
  signal L2_shift_L23_n_275, L2_shift_L23_n_276, L2_shift_L23_n_277, L2_shift_L23_n_278, L2_shift_L23_n_279 : std_logic;
  signal L2_shift_L23_n_280, L2_shift_L23_n_281, L2_shift_L23_n_282, L2_shift_L23_n_283, L2_shift_L23_n_284 : std_logic;
  signal L2_shift_L23_n_285, L2_shift_L23_n_286, L2_shift_L23_n_288, L2_shift_L23_n_289, L2_shift_L23_n_290 : std_logic;
  signal L2_shift_L23_n_291, L2_shift_L23_n_292, L2_shift_L23_n_293, L2_shift_L23_n_296, L2_shift_L23_n_297 : std_logic;
  signal L2_shift_L23_n_298, L2_shift_L23_n_299, L2_shift_L23_n_300, L2_shift_L23_n_301, L2_shift_L23_n_302 : std_logic;
  signal L2_shift_L23_n_303, L2_shift_L23_n_304, L2_shift_L23_n_305, L2_shift_L23_n_306, L2_shift_L23_n_307 : std_logic;
  signal L2_shift_L23_n_308, L2_shift_L23_n_309, L2_shift_L23_n_310, L2_shift_L23_n_311, L2_shift_L23_n_312 : std_logic;
  signal L2_shift_L23_n_313, L2_shift_L23_n_314, L2_shift_L23_n_315, L2_shift_L23_n_316, L2_shift_L23_n_317 : std_logic;
  signal L2_shift_L23_n_318, L2_shift_L23_n_319, L2_shift_L23_n_320, L2_shift_L23_n_321, L2_shift_L23_n_322 : std_logic;
  signal L2_shift_L23_n_323, L2_shift_L23_n_324, L2_shift_L23_n_325, L2_shift_L23_n_326, L2_shift_L23_n_327 : std_logic;
  signal L2_shift_L23_n_328, L2_shift_L23_n_329, L2_shift_L23_n_330, L2_shift_L23_n_331, L2_shift_L23_n_390 : std_logic;
  signal L2_shift_L23_n_394, L2_shift_L23_n_396, L2_shift_L23_n_397, L2_shift_L23_n_398, L2_shift_L23_n_399 : std_logic;
  signal L2_shift_L31_n_0, L2_shift_L31_n_1, L2_shift_L31_n_2, L2_shift_L31_n_3, L2_shift_L31_n_4 : std_logic;
  signal L2_shift_L31_n_5, L2_shift_L31_n_6, L2_shift_L31_n_7, L2_shift_L31_n_8, L2_shift_L31_n_9 : std_logic;
  signal L2_shift_L31_n_10, L2_shift_L33_n_0, L2_shift_L33_n_1, L2_shift_L33_n_2, L2_shift_L33_n_3 : std_logic;
  signal L2_shift_L33_n_4, L2_shift_L33_n_5, L2_shift_L33_n_6, L2_shift_L33_n_7, L2_shift_L33_n_8 : std_logic;
  signal L2_shift_L33_n_9, L2_shift_L33_n_10, L2_shift_L33_n_11, L2_shift_L33_n_12, L2_shift_L33_n_13 : std_logic;
  signal L2_shift_L33_n_14, L2_shift_L33_n_15, L2_shift_L33_n_16, L2_shift_L33_n_17, L2_shift_L33_n_18 : std_logic;
  signal L2_shift_L33_n_19, L2_shift_L33_n_20, L2_shift_L33_n_21, L2_shift_L33_n_22, L2_shift_L33_n_23 : std_logic;
  signal L2_shift_L33_n_24, L2_shift_L33_n_25, L2_shift_L33_n_26, L2_shift_L33_n_27, L2_shift_L33_n_28 : std_logic;
  signal L2_shift_L33_n_29, L2_shift_L33_n_30, L2_shift_L33_n_31, L2_shift_L33_n_32, L2_shift_L33_n_33 : std_logic;
  signal L2_shift_L33_n_34, L2_shift_L33_n_35, L2_shift_L33_n_36, L2_shift_L33_n_37, L2_shift_L33_n_38 : std_logic;
  signal L2_shift_L33_n_39, L2_shift_L33_n_40, L2_shift_L33_n_41, L2_shift_L33_n_42, L2_shift_L33_n_43 : std_logic;
  signal L2_shift_L33_n_44, L2_shift_L33_n_45, L2_shift_L33_n_46, L2_shift_L33_n_47, L2_shift_L33_n_48 : std_logic;
  signal L2_shift_L33_n_49, L2_shift_L33_n_50, L2_shift_L33_n_51, L2_shift_L33_n_52, L2_shift_L33_n_53 : std_logic;
  signal L2_shift_L33_n_54, L2_shift_L33_n_55, L2_shift_L33_n_56, L2_shift_L33_n_57, L2_shift_L33_n_58 : std_logic;
  signal L2_shift_L33_n_59, L2_shift_L33_n_61, L2_shift_L33_n_62, L2_shift_L33_n_63, L2_shift_L33_n_64 : std_logic;
  signal L2_shift_L33_n_65, L2_shift_L33_n_66, L2_shift_L33_n_67, L2_shift_L33_n_68, L2_shift_L33_n_69 : std_logic;
  signal L2_shift_L33_n_70, L2_shift_L33_n_71, L2_shift_L33_n_72, L2_shift_L33_n_73, L2_shift_L33_n_74 : std_logic;
  signal L2_shift_L33_n_75, L2_shift_L33_n_76, L2_shift_L33_n_77, L2_shift_L33_n_78, L2_shift_L33_n_79 : std_logic;
  signal L2_shift_L33_n_80, L2_shift_L33_n_81, L2_shift_L33_n_82, L2_shift_L33_n_83, L2_shift_L33_n_84 : std_logic;
  signal L2_shift_L33_n_85, L2_shift_L33_n_86, L2_shift_L33_n_87, L2_shift_L33_n_88, L2_shift_L33_n_89 : std_logic;
  signal L2_shift_L33_n_90, L2_shift_L33_n_91, L2_shift_L33_n_92, L2_shift_L33_n_93, L2_shift_L33_n_94 : std_logic;
  signal L2_shift_L33_n_95, L2_shift_L33_n_96, L2_shift_L33_n_97, L2_shift_L33_n_98, L2_shift_L33_n_99 : std_logic;
  signal L2_shift_L33_n_100, L2_shift_L33_n_101, L2_shift_L33_n_102, L2_shift_L33_n_103, L2_shift_L33_n_104 : std_logic;
  signal L2_shift_L33_n_105, L2_shift_L33_n_106, L2_shift_L33_n_107, L2_shift_L33_n_108, L2_shift_L33_n_109 : std_logic;
  signal L2_shift_L33_n_110, L2_shift_L33_n_111, L2_shift_L33_n_112, L2_shift_L33_n_113, L2_shift_L33_n_114 : std_logic;
  signal L2_shift_L33_n_115, L2_shift_L33_n_116, L2_shift_L33_n_117, L2_shift_L33_n_118, L2_shift_L33_n_119 : std_logic;
  signal L2_shift_L33_n_120, L2_shift_L33_n_121, L2_shift_L33_n_122, L2_shift_L33_n_123, L2_shift_L33_n_124 : std_logic;
  signal L2_shift_L33_n_125, L2_shift_L33_n_126, L2_shift_L33_n_127, L2_shift_L33_n_128, L2_shift_L33_n_129 : std_logic;
  signal L2_shift_L33_n_131, L2_shift_L33_n_132, L2_shift_L33_n_133, L2_shift_L33_n_134, L2_shift_L33_n_135 : std_logic;
  signal L2_shift_L33_n_136, L2_shift_L33_n_137, L2_shift_L33_n_138, L2_shift_L33_n_139, L2_shift_L33_n_140 : std_logic;
  signal L2_shift_L33_n_141, L2_shift_L33_n_142, L2_shift_L33_n_143, L2_shift_L33_n_144, L2_shift_L33_n_145 : std_logic;
  signal L2_shift_L33_n_146, L2_shift_L33_n_147, L2_shift_L33_n_149, L2_shift_L33_n_150, L2_shift_L33_n_151 : std_logic;
  signal L2_shift_L33_n_152, L2_shift_L33_n_153, L2_shift_L33_n_154, L2_shift_L33_n_155, L2_shift_L33_n_156 : std_logic;
  signal L2_shift_L33_n_157, L2_shift_L33_n_159, L2_shift_L33_n_160, L2_shift_L33_n_161, L2_shift_L33_n_162 : std_logic;
  signal L2_shift_L33_n_163, L2_shift_L33_n_164, L2_shift_L33_n_165, L2_shift_L33_n_166, L2_shift_L33_n_167 : std_logic;
  signal L2_shift_L33_n_168, L2_shift_L33_n_169, L2_shift_L33_n_170, L2_shift_L33_n_171, L2_shift_L33_n_172 : std_logic;
  signal L2_shift_L33_n_173, L2_shift_L33_n_174, L2_shift_L33_n_175, L2_shift_L33_n_176, L2_shift_L33_n_177 : std_logic;
  signal L2_shift_L33_n_178, L2_shift_L33_n_179, L2_shift_L33_n_180, L2_shift_L33_n_181, L2_shift_L33_n_182 : std_logic;
  signal L2_shift_L33_n_183, L2_shift_L33_n_184, L2_shift_L33_n_185, L2_shift_L33_n_186, L2_shift_L33_n_187 : std_logic;
  signal L2_shift_L33_n_188, L2_shift_L33_n_189, L2_shift_L33_n_190, L2_shift_L33_n_191, L2_shift_L33_n_192 : std_logic;
  signal L2_shift_L33_n_193, L2_shift_L33_n_194, L2_shift_L33_n_195, L2_shift_L33_n_196, L2_shift_L33_n_197 : std_logic;
  signal L2_shift_L33_n_198, L2_shift_L33_n_199, L2_shift_L33_n_200, L2_shift_L33_n_201, L2_shift_L33_n_202 : std_logic;
  signal L2_shift_L33_n_203, L2_shift_L33_n_204, L2_shift_L33_n_205, L2_shift_L33_n_206, L2_shift_L33_n_207 : std_logic;
  signal L2_shift_L33_n_208, L2_shift_L33_n_209, L2_shift_L33_n_210, L2_shift_L33_n_211, L2_shift_L33_n_212 : std_logic;
  signal L2_shift_L33_n_213, L2_shift_L33_n_214, L2_shift_L33_n_215, L2_shift_L33_n_216, L2_shift_L33_n_217 : std_logic;
  signal L2_shift_L33_n_218, L2_shift_L33_n_219, L2_shift_L33_n_220, L2_shift_L33_n_221, L2_shift_L33_n_222 : std_logic;
  signal L2_shift_L33_n_223, L2_shift_L33_n_224, L2_shift_L33_n_225, L2_shift_L33_n_226, L2_shift_L33_n_227 : std_logic;
  signal L2_shift_L33_n_228, L2_shift_L33_n_229, L2_shift_L33_n_230, L2_shift_L33_n_231, L2_shift_L33_n_232 : std_logic;
  signal L2_shift_L33_n_233, L2_shift_L33_n_235, L2_shift_L33_n_236, L2_shift_L33_n_237, L2_shift_L33_n_238 : std_logic;
  signal L2_shift_L33_n_239, L2_shift_L33_n_240, L2_shift_L33_n_241, L2_shift_L33_n_242, L2_shift_L33_n_243 : std_logic;
  signal L2_shift_L33_n_244, L2_shift_L33_n_245, L2_shift_L33_n_246, L2_shift_L33_n_247, L2_shift_L33_n_248 : std_logic;
  signal L2_shift_L33_n_249, L2_shift_L33_n_250, L2_shift_L33_n_251, L2_shift_L33_n_252, L2_shift_L33_n_253 : std_logic;
  signal L2_shift_L33_n_254, L2_shift_L33_n_255, L2_shift_L33_n_256, L2_shift_L33_n_257, L2_shift_L33_n_258 : std_logic;
  signal L2_shift_L33_n_259, L2_shift_L33_n_260, L2_shift_L33_n_261, L2_shift_L33_n_262, L2_shift_L33_n_263 : std_logic;
  signal L2_shift_L33_n_264, L2_shift_L33_n_265, L2_shift_L33_n_266, L2_shift_L33_n_267, L2_shift_L33_n_268 : std_logic;
  signal L2_shift_L33_n_269, L2_shift_L33_n_270, L2_shift_L33_n_271, L2_shift_L33_n_272, L2_shift_L33_n_273 : std_logic;
  signal L2_shift_L33_n_274, L2_shift_L33_n_275, L2_shift_L33_n_276, L2_shift_L33_n_277, L2_shift_L33_n_278 : std_logic;
  signal L2_shift_L33_n_279, L2_shift_L33_n_280, L2_shift_L33_n_281, L2_shift_L33_n_282, L2_shift_L33_n_283 : std_logic;
  signal L2_shift_L33_n_285, L2_shift_L33_n_286, L2_shift_L33_n_287, L2_shift_L33_n_288, L2_shift_L33_n_289 : std_logic;
  signal L2_shift_L33_n_290, L2_shift_L33_n_293, L2_shift_L33_n_294, L2_shift_L33_n_295, L2_shift_L33_n_296 : std_logic;
  signal L2_shift_L33_n_297, L2_shift_L33_n_298, L2_shift_L33_n_299, L2_shift_L33_n_300, L2_shift_L33_n_301 : std_logic;
  signal L2_shift_L33_n_302, L2_shift_L33_n_303, L2_shift_L33_n_304, L2_shift_L33_n_305, L2_shift_L33_n_306 : std_logic;
  signal L2_shift_L33_n_307, L2_shift_L33_n_308, L2_shift_L33_n_309, L2_shift_L33_n_310, L2_shift_L33_n_311 : std_logic;
  signal L2_shift_L33_n_312, L2_shift_L33_n_313, L2_shift_L33_n_314, L2_shift_L33_n_315, L2_shift_L33_n_316 : std_logic;
  signal L2_shift_L33_n_317, L2_shift_L33_n_318, L2_shift_L33_n_319, L2_shift_L33_n_320, L2_shift_L33_n_321 : std_logic;
  signal L2_shift_L33_n_322, L2_shift_L33_n_323, L2_shift_L33_n_324, L2_shift_L33_n_325, L2_shift_L33_n_326 : std_logic;
  signal L2_shift_L33_n_327, L2_shift_L33_n_328, L2_shift_L33_n_387, L2_shift_L33_n_391, L2_shift_L33_n_393 : std_logic;
  signal L2_shift_L33_n_394, L2_shift_L33_n_395, L2_shift_L33_n_396, L2_shift_gg_pos_load, L2_shift_gg_pos_reset : std_logic;
  signal L2_shift_gr_pos_load, L2_shift_gr_pos_reset, L2_shift_pacman_pos_load, L2_shift_pacman_pos_reset, L2_shift_shift_clock_reset : std_logic;
  signal L2_shift_shift_clock_reset_gg, L2_shift_shift_clock_reset_gr, L2_shift_shift_pulse, L2_shift_shift_pulse_gg, L2_shift_shift_pulse_gr : std_logic;
  signal L2_user_reset_new, L2_vidcontrol_n_3, L2_vidcontrol_n_4, L2_vidcontrol_n_5, L2_vidcontrol_n_6 : std_logic;
  signal L2_vidcontrol_n_7, L2_vidcontrol_n_8, L2_vidcontrol_n_9, L2_vidcontrol_n_10, L2_vidcontrol_n_11 : std_logic;
  signal L2_vidcontrol_n_12, L2_vidcontrol_n_13, L2_vidcontrol_n_14, L2_vidcontrol_n_15, L2_vidcontrol_n_16 : std_logic;
  signal L2_vidcontrol_n_18, L2_vidcontrol_n_19, L2_vidcontrol_n_20, L2_vidcontrol_n_21, L2_vidcontrol_n_22 : std_logic;
  signal L2_vidcontrol_n_23, L2_vidcontrol_n_24, L2_vidcontrol_n_25, L2_vidcontrol_n_26, L2_vidcontrol_n_27 : std_logic;
  signal L2_vidcontrol_n_28, L2_vidcontrol_n_29, L2_vidcontrol_n_30, L2_vidcontrol_n_31, L2_vidcontrol_n_32 : std_logic;
  signal L2_vidcontrol_n_33, L2_vidcontrol_n_34, L2_vidcontrol_n_35, L2_vidcontrol_n_36, L2_vidcontrol_n_37 : std_logic;
  signal L2_vidcontrol_n_38, L2_vidcontrol_n_39, L2_vidcontrol_n_40, L2_vidcontrol_n_41, L2_vidcontrol_n_42 : std_logic;
  signal L2_vidcontrol_n_43, L2_vidcontrol_n_44, L2_vidcontrol_n_45, L2_vidcontrol_n_46, L2_vidcontrol_n_47 : std_logic;
  signal L2_vidcontrol_n_49, L2_vidcontrol_n_50, L2_vidcontrol_n_51, L2_vidcontrol_n_52, L2_vidcontrol_n_53 : std_logic;
  signal L2_vidcontrol_n_54, L2_vidcontrol_n_55, L2_vidcontrol_n_56, L2_vidcontrol_n_57, L2_vidcontrol_n_58 : std_logic;
  signal L2_vidcontrol_n_59, L2_vidcontrol_n_60, L2_vidcontrol_n_72, L2_vidcontrol_n_76, L2_vidcontrol_n_77 : std_logic;
  signal L2_vidcontrol_n_78, L2_vidcontrol_n_79, L2_vidcontrol_n_82, L2_vidcontrol_n_83, L2_vidcontrol_n_123 : std_logic;
  signal L2_vidcontrol_n_124, L2_vidcontrol_n_125, L2_vidcontrol_n_126, UNCONNECTED, UNCONNECTED0 : std_logic;
  signal UNCONNECTED1, UNCONNECTED2, calc_start_game_int, game_over_out_int, score_pulse_int : std_logic;

begin

  L1_g1280 : INVD1BWP7T port map(I => calc_start_game_int, ZN => L1_n_23);
  L1_g4970 : AO31D1BWP7T port map(A1 => L1_coin_present, A2 => L1_n_106, A3 => L1_n_96, B => L1_pos_is_wall, Z => cell_type_int(2));
  L1_g4971 : AOI21D0BWP7T port map(A1 => L1_n_110, A2 => L1_n_96, B => L1_pos_is_wall, ZN => cell_type_int(0));
  L1_g4972 : AO21D0BWP7T port map(A1 => L1_n_105, A2 => L1_n_96, B => L1_pos_is_wall, Z => cell_type_int(1));
  L1_g4973 : IND4D0BWP7T port map(A1 => L1_n_175, B1 => L1_n_173, B2 => L1_n_177, B3 => L1_n_178, ZN => L1_pos_is_wall);
  L1_g4974 : AOI31D0BWP7T port map(A1 => L1_n_163, A2 => L1_n_118, A3 => L1_n_123, B => L1_n_176, ZN => L1_n_178);
  L1_g4975 : AOI31D0BWP7T port map(A1 => L1_n_171, A2 => L1_n_136, A3 => L1_n_131, B => L1_n_164, ZN => L1_n_177);
  L1_g4976 : OAI221D0BWP7T port map(A1 => L1_n_167, A2 => L1_n_125, B1 => L1_n_143, B2 => L1_n_158, C => L1_n_174, ZN => L1_n_176);
  L1_g4977 : OAI32D1BWP7T port map(A1 => L1_n_130, A2 => L1_n_144, A3 => L1_n_166, B1 => L1_n_129, B2 => L1_n_169, ZN => L1_n_175);
  L1_g4978 : AOI31D0BWP7T port map(A1 => L1_n_160, A2 => L1_n_136, A3 => L1_n_129, B => L1_n_172, ZN => L1_n_174);
  L1_g4979 : OA33D0BWP7T port map(A1 => L1_n_118, A2 => L1_n_128, A3 => L1_n_165, B1 => L1_n_131, B2 => L1_n_143, B3 => L1_n_162, Z => L1_n_173);
  L1_g4980 : NR3D0BWP7T port map(A1 => L1_n_168, A2 => L1_n_144, A3 => L1_n_131, ZN => L1_n_172);
  L1_g4981 : AO21D0BWP7T port map(A1 => L1_n_129, A2 => L1_n_135, B => L1_n_170, Z => L1_n_171);
  L1_g4982 : OAI31D0BWP7T port map(A1 => L1_n_126, A2 => L1_n_140, A3 => L1_n_141, B => L1_n_168, ZN => L1_n_170);
  L1_g4983 : OAI211D1BWP7T port map(A1 => L1_n_152, A2 => L1_n_161, B => L1_n_136, C => L1_n_130, ZN => L1_n_169);
  L1_g4984 : ND4D0BWP7T port map(A1 => L1_n_154, A2 => L1_n_118, A3 => L1_n_119, A4 => L1_n_123, ZN => L1_n_167);
  L1_g4985 : NR3D0BWP7T port map(A1 => L1_n_159, A2 => L1_n_156, A3 => L1_n_151, ZN => L1_n_168);
  L1_g4986 : AOI211XD0BWP7T port map(A1 => L1_n_149, A2 => L1_n_141, B => L1_n_161, C => L1_n_155, ZN => L1_n_166);
  L1_g4987 : AOI22D0BWP7T port map(A1 => L1_n_159, A2 => L1_n_141, B1 => L1_n_149, B2 => L1_n_147, ZN => L1_n_165);
  L1_g4988 : INR4D0BWP7T port map(A1 => L1_n_119, B1 => L1_n_118, B2 => L1_n_125, B3 => L1_n_150, ZN => L1_n_164);
  L1_g4989 : NR2D1BWP7T port map(A1 => L1_n_157, A2 => L1_n_128, ZN => L1_n_163);
  L1_g4990 : AOI211XD0BWP7T port map(A1 => L1_n_153, A2 => L1_n_140, B => L1_n_156, C => L1_n_152, ZN => L1_n_162);
  L1_g4991 : AO21D0BWP7T port map(A1 => L1_n_149, A2 => L1_n_140, B => L1_n_155, Z => L1_n_160);
  L1_g4992 : AN2D1BWP7T port map(A1 => L1_n_156, A2 => L1_n_140, Z => L1_n_161);
  L1_g4993 : AOI21D0BWP7T port map(A1 => L1_n_149, A2 => L1_n_139, B => L1_n_151, ZN => L1_n_158);
  L1_g4994 : INR3D0BWP7T port map(A1 => L1_n_150, B1 => L1_n_152, B2 => L1_n_149, ZN => L1_n_157);
  L1_g4995 : AO21D0BWP7T port map(A1 => L1_n_153, A2 => L1_n_139, B => L1_n_155, Z => L1_n_159);
  L1_g4996 : INR2D1BWP7T port map(A1 => L1_n_153, B1 => L1_n_141, ZN => L1_n_156);
  L1_g4997 : OAI22D0BWP7T port map(A1 => L1_n_148, A2 => L1_n_146, B1 => L1_n_142, B2 => L1_n_126, ZN => L1_n_154);
  L1_g4998 : NR3D0BWP7T port map(A1 => L1_n_145, A2 => L1_n_140, A3 => L1_n_126, ZN => L1_n_155);
  L1_g4999 : INR2D1BWP7T port map(A1 => L1_n_126, B1 => L1_n_146, ZN => L1_n_153);
  L1_g5000 : NR2D1BWP7T port map(A1 => L1_n_148, A2 => L1_n_126, ZN => L1_n_152);
  L1_g5001 : INR2D1BWP7T port map(A1 => L1_n_147, B1 => L1_n_126, ZN => L1_n_151);
  L1_g5002 : ND2D1BWP7T port map(A1 => L1_n_147, A2 => L1_n_145, ZN => L1_n_150);
  L1_g5003 : NR2D1BWP7T port map(A1 => L1_n_146, A2 => L1_n_126, ZN => L1_n_149);
  L1_g5004 : NR2XD0BWP7T port map(A1 => L1_n_141, A2 => L1_n_139, ZN => L1_n_148);
  L1_g5005 : INVD0BWP7T port map(I => L1_n_146, ZN => L1_n_145);
  L1_g5006 : NR2D1BWP7T port map(A1 => L1_n_142, A2 => L1_n_139, ZN => L1_n_147);
  L1_g5007 : OAI211D1BWP7T port map(A1 => L1_n_120, A2 => L1_n_134, B => L1_n_138, C => L1_n_135, ZN => L1_n_146);
  L1_g5008 : ND2D1BWP7T port map(A1 => L1_n_137, A2 => L1_n_129, ZN => L1_n_144);
  L1_g5009 : IND2D1BWP7T port map(A1 => L1_n_129, B1 => L1_n_137, ZN => L1_n_143);
  L1_g5010 : INVD1BWP7T port map(I => L1_n_142, ZN => L1_n_141);
  L1_g5011 : INVD1BWP7T port map(I => L1_n_140, ZN => L1_n_139);
  L1_g5012 : CKXOR2D1BWP7T port map(A1 => L1_n_134, A2 => L1_n_109, Z => L1_n_142);
  L1_g5013 : MAOI22D0BWP7T port map(A1 => L1_n_134, A2 => L1_n_111, B1 => L1_n_134, B2 => L1_n_111, ZN => L1_n_140);
  L1_g5014 : ND2D1BWP7T port map(A1 => L1_n_134, A2 => L1_n_120, ZN => L1_n_138);
  L1_g5015 : NR2D1BWP7T port map(A1 => L1_n_132, A2 => L1_n_123, ZN => L1_n_137);
  L1_g5016 : NR2D1BWP7T port map(A1 => L1_n_133, A2 => L1_n_123, ZN => L1_n_136);
  L1_g5017 : ND2D1BWP7T port map(A1 => L1_n_127, A2 => L1_n_126, ZN => L1_n_135);
  L1_g5018 : AOI21D0BWP7T port map(A1 => L1_n_126, A2 => L1_n_120, B => L1_n_127, ZN => L1_n_134);
  L1_g5019 : INVD0BWP7T port map(I => L1_n_132, ZN => L1_n_133);
  L1_g5020 : INVD0BWP7T port map(I => L1_n_131, ZN => L1_n_130);
  L1_g5021 : MAOI22D0BWP7T port map(A1 => L1_n_125, A2 => L1_n_117, B1 => L1_n_125, B2 => L1_n_117, ZN => L1_n_132);
  L1_g5022 : MOAI22D0BWP7T port map(A1 => L1_n_125, A2 => L1_n_107, B1 => L1_n_125, B2 => L1_n_107, ZN => L1_n_131);
  L1_g5023 : MOAI22D0BWP7T port map(A1 => L1_n_125, A2 => L1_n_108, B1 => L1_n_125, B2 => L1_n_108, ZN => L1_n_129);
  L1_g5024 : OR2D1BWP7T port map(A1 => L1_n_125, A2 => L1_n_119, Z => L1_n_128);
  L1_g5025 : AO221D0BWP7T port map(A1 => L1_row_new_pacman(4), A2 => L1_n_35, B1 => ycoordinates_int(4), B2 => L1_n_23, C => L1_n_124, Z => L1_n_127);
  L1_g5026 : ND3D0BWP7T port map(A1 => L1_n_90, A2 => L1_n_121, A3 => L1_n_38, ZN => L1_n_126);
  L1_g5027 : AO22D0BWP7T port map(A1 => L1_n_190, A2 => L1_n_83, B1 => L1_n_82, B2 => L1_row_old_ghost1(4), Z => L1_n_124);
  L1_g5028 : AO222D0BWP7T port map(A1 => L1_col_new_pacman(4), A2 => L1_n_35, B1 => L1_n_184, B2 => L1_n_31, C1 => xcoordinates_int(4), C2 => L1_n_23, Z => L1_n_125);
  L1_g5029 : ND2D1BWP7T port map(A1 => L1_n_122, A2 => L1_n_38, ZN => L1_n_123);
  L1_g5030 : AOI222D0BWP7T port map(A1 => L1_n_35, A2 => L1_col_new_pacman(3), B1 => xcoordinates_int(3), B2 => L1_n_23, C1 => L1_n_31, C2 => L1_n_186, ZN => L1_n_122);
  L1_g5031 : OAI222D0BWP7T port map(A1 => L1_n_114, A2 => L1_n_37, B1 => L1_n_36, B2 => L1_n_115, C1 => L1_n_61, C2 => L1_n_15, ZN => L1_n_190);
  L1_g5032 : AOI22D0BWP7T port map(A1 => L1_n_185, A2 => L1_n_83, B1 => ycoordinates_int(3), B2 => L1_n_23, ZN => L1_n_121);
  L1_g5033 : OAI222D0BWP7T port map(A1 => L1_n_114, A2 => L1_n_86, B1 => L1_n_88, B2 => L1_n_115, C1 => L1_n_81, C2 => L1_n_20, ZN => L1_n_184);
  L1_g5034 : ND3D0BWP7T port map(A1 => L1_n_89, A2 => L1_n_116, A3 => L1_n_38, ZN => L1_n_120);
  L1_g5035 : CKXOR2D1BWP7T port map(A1 => L1_n_117, A2 => L1_n_108, Z => L1_n_119);
  L1_g5036 : XNR2D1BWP7T port map(A1 => L1_n_117, A2 => L1_n_107, ZN => L1_n_118);
  L1_g5037 : OAI222D0BWP7T port map(A1 => L1_n_113, A2 => L1_n_37, B1 => L1_n_36, B2 => L1_n_103, C1 => L1_n_61, C2 => L1_n_16, ZN => L1_n_185);
  L1_g5038 : OAI222D0BWP7T port map(A1 => L1_n_113, A2 => L1_n_86, B1 => L1_n_88, B2 => L1_n_103, C1 => L1_n_81, C2 => L1_n_29, ZN => L1_n_186);
  L1_g5039 : AOI22D0BWP7T port map(A1 => L1_n_181, A2 => L1_n_83, B1 => ycoordinates_int(2), B2 => L1_n_23, ZN => L1_n_116);
  L1_g5040 : AOI222D0BWP7T port map(A1 => L1_n_31, A2 => L1_n_187, B1 => L1_n_35, B2 => L1_col_new_pacman(2), C1 => xcoordinates_int(2), C2 => L1_n_23, ZN => L1_n_117);
  L1_g5041 : MAOI22D0BWP7T port map(A1 => L1_n_100, A2 => L1_n_69, B1 => L1_n_100, B2 => L1_n_69, ZN => L1_n_115);
  L1_g5042 : MAOI22D0BWP7T port map(A1 => L1_n_112, A2 => L1_n_70, B1 => L1_n_112, B2 => L1_n_70, ZN => L1_n_114);
  L1_g5043 : HA1D0BWP7T port map(A => L1_n_55, B => L1_n_92, CO => L1_n_112, S => L1_n_113);
  L1_g5044 : OAI21D0BWP7T port map(A1 => L1_coin_present, A2 => L1_n_99, B => L1_n_97, ZN => L1_n_110);
  L1_g5045 : AO221D0BWP7T port map(A1 => L1_n_35, A2 => L1_row_new_pacman(1), B1 => ycoordinates_int(1), B2 => L1_n_23, C => L1_n_101, Z => L1_n_111);
  L1_g5046 : AOI222D0BWP7T port map(A1 => L1_n_21, A2 => L1_n_98, B1 => ycoordinates_int(0), B2 => L1_n_23, C1 => L1_n_66, C2 => L1_row_new_pacman(0), ZN => L1_n_109);
  L1_g5047 : OAI222D0BWP7T port map(A1 => L1_n_95, A2 => L1_n_37, B1 => L1_n_36, B2 => L1_n_94, C1 => L1_n_61, C2 => L1_n_26, ZN => L1_n_181);
  L1_g5048 : OAI222D0BWP7T port map(A1 => L1_n_95, A2 => L1_n_86, B1 => L1_n_88, B2 => L1_n_94, C1 => L1_n_81, C2 => L1_n_28, ZN => L1_n_187);
  L1_g5049 : AO221D0BWP7T port map(A1 => L1_n_66, A2 => L1_col_new_pacman(1), B1 => xcoordinates_int(1), B2 => L1_n_23, C => L1_n_104, Z => L1_n_108);
  L1_g5050 : AO221D0BWP7T port map(A1 => L1_n_66, A2 => L1_col_new_pacman(0), B1 => xcoordinates_int(0), B2 => L1_n_23, C => L1_n_102, Z => L1_n_107);
  L1_g5051 : INVD0BWP7T port map(I => L1_n_105, ZN => L1_n_106);
  L1_g5052 : AN3D0BWP7T port map(A1 => L1_n_31, A2 => L1_n_21, A3 => L1_n_188, Z => L1_n_104);
  L1_g5053 : IND2D1BWP7T port map(A1 => L1_n_99, B1 => L1_n_97, ZN => L1_n_105);
  L1_g5054 : AN3D0BWP7T port map(A1 => L1_n_31, A2 => L1_n_21, A3 => L1_n_189, Z => L1_n_102);
  L1_g5055 : AO22D0BWP7T port map(A1 => L1_n_182, A2 => L1_n_83, B1 => L1_n_82, B2 => L1_row_old_ghost1(1), Z => L1_n_101);
  L1_g5056 : MAOI22D0BWP7T port map(A1 => L1_n_93, A2 => L1_n_64, B1 => L1_n_93, B2 => L1_n_64, ZN => L1_n_103);
  L1_g5057 : INR2XD0BWP7T port map(A1 => L1_n_93, B1 => L1_n_64, ZN => L1_n_100);
  L1_g5058 : NR4D0BWP7T port map(A1 => L1_n_91, A2 => xcoordinates_int(0), A3 => L1_n_24, A4 => xcoordinates_int(1), ZN => L1_n_99);
  L1_g5059 : OAI222D0BWP7T port map(A1 => L1_n_86, A2 => L1_n_62, B1 => L1_n_60, B2 => L1_n_88, C1 => L1_n_81, C2 => L1_n_27, ZN => L1_n_189);
  L1_g5060 : OAI222D0BWP7T port map(A1 => L1_n_84, A2 => L1_n_37, B1 => L1_n_36, B2 => L1_n_80, C1 => L1_n_61, C2 => L1_n_25, ZN => L1_n_182);
  L1_g5061 : AO22D0BWP7T port map(A1 => L1_n_183, A2 => L1_n_83, B1 => L1_n_82, B2 => L1_row_old_ghost1(0), Z => L1_n_98);
  L1_g5062 : OAI222D0BWP7T port map(A1 => L1_n_84, A2 => L1_n_86, B1 => L1_n_88, B2 => L1_n_80, C1 => L1_n_81, C2 => L1_n_19, ZN => L1_n_188);
  L1_g5063 : OAI211D1BWP7T port map(A1 => L1_col_old_ghost1(2), A2 => L1_n_24, B => L1_n_85, C => L1_n_78, ZN => L1_n_97);
  L1_g5064 : ND4D0BWP7T port map(A1 => L1_n_76, A2 => L1_n_77, A3 => L1_n_72, A4 => L1_n_54, ZN => L1_n_96);
  L1_g5065 : AOI21D0BWP7T port map(A1 => L1_n_74, A2 => L1_n_68, B => L1_n_92, ZN => L1_n_95);
  L1_g5066 : MAOI22D0BWP7T port map(A1 => L1_n_73, A2 => L1_n_65, B1 => L1_n_73, B2 => L1_n_65, ZN => L1_n_94);
  L1_g5067 : ND2D1BWP7T port map(A1 => L1_n_87, A2 => xcoordinates_int(3), ZN => L1_n_91);
  L1_g5068 : INR2XD0BWP7T port map(A1 => L1_n_73, B1 => L1_n_65, ZN => L1_n_93);
  L1_g5069 : NR2XD0BWP7T port map(A1 => L1_n_74, A2 => L1_n_68, ZN => L1_n_92);
  L1_g5070 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(3), A2 => L1_n_82, B1 => L1_n_35, B2 => L1_row_new_pacman(3), ZN => L1_n_90);
  L1_g5071 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(2), A2 => L1_n_82, B1 => L1_n_35, B2 => L1_row_new_pacman(2), ZN => L1_n_89);
  L1_g5072 : OAI222D0BWP7T port map(A1 => L1_n_62, A2 => L1_n_37, B1 => L1_n_36, B2 => L1_n_60, C1 => L1_n_61, C2 => L1_n_18, ZN => L1_n_183);
  L1_g5073 : NR4D0BWP7T port map(A1 => L1_n_57, A2 => ycoordinates_int(1), A3 => ycoordinates_int(0), A4 => xcoordinates_int(4), ZN => L1_n_87);
  L1_g5074 : ND3D0BWP7T port map(A1 => L1_n_32, A2 => L1_n_22, A3 => L1_L3a_move(0), ZN => L1_n_88);
  L1_g5075 : AOI211XD0BWP7T port map(A1 => L1_n_24, A2 => L1_col_old_ghost1(2), B => L1_n_79, C => L1_n_48, ZN => L1_n_85);
  L1_g5076 : IND3D0BWP7T port map(A1 => L1_L3a_move(0), B1 => L1_L3a_move(2), B2 => L1_n_32, ZN => L1_n_86);
  L1_g5077 : OA21D0BWP7T port map(A1 => L1_n_63, A2 => L1_n_71, B => L1_n_74, Z => L1_n_84);
  L1_g5078 : AN2D1BWP7T port map(A1 => L1_n_31, A2 => L1_n_33, Z => L1_n_83);
  L1_g5079 : INR2D1BWP7T port map(A1 => L1_n_31, B1 => L1_n_33, ZN => L1_n_82);
  L1_g5080 : AOI211D0BWP7T port map(A1 => L1_L3a_move(2), A2 => L1_L3a_move(0), B => L1_n_33, C => L1_n_75, ZN => L1_n_81);
  L1_g5081 : ND4D0BWP7T port map(A1 => L1_n_40, A2 => L1_n_49, A3 => L1_n_58, A4 => L1_n_42, ZN => L1_n_79);
  L1_g5082 : NR4D0BWP7T port map(A1 => L1_n_39, A2 => L1_n_50, A3 => L1_n_51, A4 => L1_n_46, ZN => L1_n_78);
  L1_g5083 : NR3D0BWP7T port map(A1 => L1_n_41, A2 => L1_n_45, A3 => L1_n_47, ZN => L1_n_77);
  L1_g5084 : NR4D0BWP7T port map(A1 => L1_n_43, A2 => L1_n_53, A3 => L1_n_52, A4 => L1_n_56, ZN => L1_n_76);
  L1_g5085 : MAOI22D0BWP7T port map(A1 => L1_n_67, A2 => L1_n_60, B1 => L1_n_67, B2 => L1_n_60, ZN => L1_n_80);
  L1_g5086 : INVD0BWP7T port map(I => L1_n_32, ZN => L1_n_75);
  L1_g5087 : ND2D1BWP7T port map(A1 => L1_n_71, A2 => L1_n_63, ZN => L1_n_74);
  L1_g5088 : AOI211XD0BWP7T port map(A1 => L1_n_17, A2 => L1_row_old_pacman(1), B => L1_n_30, C => L1_n_44, ZN => L1_n_72);
  L1_g5089 : NR2XD0BWP7T port map(A1 => L1_n_59, A2 => L1_n_67, ZN => L1_n_73);
  L1_g5090 : INVD0BWP7T port map(I => L1_n_63, ZN => L1_n_62);
  L1_g5091 : INVD1BWP7T port map(I => L1_n_59, ZN => L1_n_60);
  L1_g5092 : MAOI22D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L1_n_29, B1 => xcoordinates_int(3), B2 => L1_n_29, ZN => L1_n_58);
  L1_g5093 : OR2D1BWP7T port map(A1 => L1_zero_coins, A2 => game_over_out_int, Z => L1_L5_n_14);
  L1_g5094 : IND3D1BWP7T port map(A1 => ycoordinates_int(4), B1 => ycoordinates_int(2), B2 => ycoordinates_int(3), ZN => L1_n_57);
  L1_g5095 : MOAI22D0BWP7T port map(A1 => L1_n_24, A2 => L1_col_old_pacman(2), B1 => L1_n_24, B2 => L1_col_old_pacman(2), ZN => L1_n_56);
  L1_g5096 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(1), A2 => L1_n_22, B1 => L1_col_old_ghost1(1), B2 => L1_L3a_move(2), ZN => L1_n_71);
  L1_g5097 : OAI22D0BWP7T port map(A1 => L1_row_old_ghost1(4), A2 => L1_L3a_move(2), B1 => L1_col_old_ghost1(4), B2 => L1_n_22, ZN => L1_n_70);
  L1_g5098 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(4), A2 => L1_L3a_move(3), B1 => L1_col_old_ghost1(4), B2 => L1_L3a_move(0), ZN => L1_n_69);
  L1_g5099 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(3), A2 => L1_n_22, B1 => L1_col_old_ghost1(3), B2 => L1_L3a_move(2), ZN => L1_n_55);
  L1_g5100 : OAI22D0BWP7T port map(A1 => L1_n_26, A2 => L1_L3a_move(2), B1 => L1_n_28, B2 => L1_n_22, ZN => L1_n_68);
  L1_g5101 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(1), A2 => L1_L3a_move(3), B1 => L1_col_old_ghost1(1), B2 => L1_L3a_move(0), ZN => L1_n_67);
  L1_g5102 : NR2D1BWP7T port map(A1 => L1_n_34, A2 => L1_ghost2_map_select, ZN => L1_n_66);
  L1_g5103 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(2), A2 => L1_L3a_move(3), B1 => L1_col_old_ghost1(2), B2 => L1_L3a_move(0), ZN => L1_n_65);
  L1_g5104 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(3), A2 => L1_L3a_move(3), B1 => L1_col_old_ghost1(3), B2 => L1_L3a_move(0), ZN => L1_n_64);
  L1_g5105 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(0), A2 => L1_n_22, B1 => L1_col_old_ghost1(0), B2 => L1_L3a_move(2), ZN => L1_n_63);
  L1_g5106 : AOI21D0BWP7T port map(A1 => L1_L3a_move(3), A2 => L1_L3a_move(1), B => L1_n_32, ZN => L1_n_61);
  L1_g5107 : AOI22D0BWP7T port map(A1 => L1_row_old_ghost1(0), A2 => L1_L3a_move(3), B1 => L1_col_old_ghost1(0), B2 => L1_L3a_move(0), ZN => L1_n_59);
  L1_g5108 : XNR2D1BWP7T port map(A1 => xcoordinates_int(1), A2 => L1_col_old_pacman(1), ZN => L1_n_54);
  L1_g5109 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(0), A2 => L1_row_old_pacman(0), Z => L1_n_53);
  L1_g5110 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(3), A2 => L1_row_old_pacman(3), Z => L1_n_52);
  L1_g5111 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L1_n_16, B1 => ycoordinates_int(3), B2 => L1_n_16, ZN => L1_n_51);
  L1_g5112 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(0), A2 => L1_n_18, B1 => ycoordinates_int(0), B2 => L1_n_18, ZN => L1_n_50);
  L1_g5113 : MAOI22D0BWP7T port map(A1 => xcoordinates_int(4), A2 => L1_n_20, B1 => xcoordinates_int(4), B2 => L1_n_20, ZN => L1_n_49);
  L1_g5114 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(2), A2 => L1_n_26, B1 => ycoordinates_int(2), B2 => L1_n_26, ZN => L1_n_48);
  L1_g5115 : CKXOR2D1BWP7T port map(A1 => xcoordinates_int(3), A2 => L1_col_old_pacman(3), Z => L1_n_47);
  L1_g5116 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(1), A2 => L1_n_19, B1 => xcoordinates_int(1), B2 => L1_n_19, ZN => L1_n_46);
  L1_g5117 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(4), A2 => L1_row_old_pacman(4), Z => L1_n_45);
  L1_g5118 : CKXOR2D1BWP7T port map(A1 => xcoordinates_int(4), A2 => L1_col_old_pacman(4), Z => L1_n_44);
  L1_g5119 : CKXOR2D1BWP7T port map(A1 => xcoordinates_int(0), A2 => L1_col_old_pacman(0), Z => L1_n_43);
  L1_g5120 : MAOI22D0BWP7T port map(A1 => ycoordinates_int(4), A2 => L1_n_15, B1 => ycoordinates_int(4), B2 => L1_n_15, ZN => L1_n_42);
  L1_g5121 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(2), A2 => L1_row_old_pacman(2), Z => L1_n_41);
  L1_g5122 : AOI22D0BWP7T port map(A1 => ycoordinates_int(1), A2 => L1_n_25, B1 => L1_n_17, B2 => L1_row_old_ghost1(1), ZN => L1_n_40);
  L1_g5123 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(0), A2 => L1_n_27, B1 => xcoordinates_int(0), B2 => L1_n_27, ZN => L1_n_39);
  L1_g5124 : INVD1BWP7T port map(I => L1_n_34, ZN => L1_n_35);
  L1_g5125 : ND2D1BWP7T port map(A1 => L1_ghost2_map_select, A2 => calc_start_game_int, ZN => L1_n_38);
  L1_g5126 : IND2D0BWP7T port map(A1 => L1_L3a_move(3), B1 => L1_L3a_move(1), ZN => L1_n_37);
  L1_g5127 : IND2D0BWP7T port map(A1 => L1_L3a_move(1), B1 => L1_L3a_move(3), ZN => L1_n_36);
  L1_g5128 : ND2D1BWP7T port map(A1 => L1_pacman_map_select, A2 => calc_start_game_int, ZN => L1_n_34);
  L1_g5129 : NR2D0BWP7T port map(A1 => L1_n_17, A2 => L1_row_old_pacman(1), ZN => L1_n_30);
  L1_g5130 : OR2D1BWP7T port map(A1 => L1_pacman_dead, A2 => reset, Z => game_over_out_int);
  L1_g5131 : NR2D0BWP7T port map(A1 => L1_L3a_move(2), A2 => L1_L3a_move(0), ZN => L1_n_33);
  L1_g5132 : NR2D0BWP7T port map(A1 => L1_L3a_move(3), A2 => L1_L3a_move(1), ZN => L1_n_32);
  L1_g5133 : NR2D1BWP7T port map(A1 => L1_pacman_map_select, A2 => L1_n_23, ZN => L1_n_31);
  L1_g5139 : INVD1BWP7T port map(I => xcoordinates_int(2), ZN => L1_n_24);
  L1_g5141 : INVD1BWP7T port map(I => L1_L3a_move(2), ZN => L1_n_22);
  L1_g5142 : INVD0BWP7T port map(I => L1_ghost2_map_select, ZN => L1_n_21);
  L1_g5146 : INVD0BWP7T port map(I => ycoordinates_int(1), ZN => L1_n_17);
  L1_L3a_L5_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L1_n_7, Q => L1_L3a_L5_state(0));
  L1_g1607 : AO221D0BWP7T port map(A1 => L1_n_185, A2 => L1_n_5, B1 => L1_row_old_ghost1(3), B2 => L1_n_4, C => game_over_out_int, Z => L1_n_13);
  L1_g1608 : AO221D0BWP7T port map(A1 => L1_n_182, A2 => L1_n_5, B1 => L1_row_old_ghost1(1), B2 => L1_n_4, C => game_over_out_int, Z => L1_n_12);
  L1_g1609 : AO221D0BWP7T port map(A1 => L1_n_183, A2 => L1_n_5, B1 => L1_row_old_ghost1(0), B2 => L1_n_4, C => game_over_out_int, Z => L1_n_11);
  L1_g1612 : AO221D0BWP7T port map(A1 => L1_n_1, A2 => L1_n_188, B1 => L1_n_2, B2 => L1_col_old_ghost1(1), C => game_over_out_int, Z => L1_n_10);
  L1_g1613 : AO221D0BWP7T port map(A1 => L1_n_1, A2 => L1_n_189, B1 => L1_n_2, B2 => L1_col_old_ghost1(0), C => game_over_out_int, Z => L1_n_9);
  L1_g1614 : AO221D0BWP7T port map(A1 => L1_n_186, A2 => L1_n_1, B1 => L1_n_2, B2 => L1_col_old_ghost1(3), C => game_over_out_int, Z => L1_n_8);
  L1_g1615 : AO21D0BWP7T port map(A1 => L1_pos_is_wall, A2 => L1_n_3, B => L1_n_6, Z => L1_n_7);
  L1_L3a_L5_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => L1_n_3, Q => L1_ghost1_ready);
  L1_g1617 : INR4D0BWP7T port map(A1 => L1_ghost1_start, B1 => L1_ghost1_ready, B2 => L1_L3a_L5_state(0), B3 => game_over_out_int, ZN => L1_n_6);
  L1_g1618 : INVD1BWP7T port map(I => L1_n_5, ZN => L1_n_4);
  L1_g1619 : NR3D0BWP7T port map(A1 => L1_n_2, A2 => L1_L3a_move(0), A3 => L1_L3a_move(2), ZN => L1_n_5);
  L1_g1620 : INR3D0BWP7T port map(A1 => L1_L3a_L5_state(0), B1 => L1_ghost1_ready, B2 => game_over_out_int, ZN => L1_n_3);
  L1_g1621 : INVD1BWP7T port map(I => L1_n_2, ZN => L1_n_1);
  L1_g1622 : IND2D1BWP7T port map(A1 => L1_L3a_L5_state(0), B1 => L1_ghost1_ready, ZN => L1_n_2);
  L1_g1623 : INVD1BWP7T port map(I => game_over_out_int, ZN => L1_n_0);
  L1_L3a_L4_column_number_out_reg_3 : DFD1BWP7T port map(CP => clk, D => L1_n_8, Q => L1_col_old_ghost1(3), QN => L1_n_29);
  L1_L3a_L4_column_number_out_reg_2 : EDFKCND1BWP7T port map(CP => clk, CN => L1_n_0, D => L1_n_187, E => L1_n_1, Q => L1_col_old_ghost1(2), QN => L1_n_28);
  L1_L3a_L4_column_number_out_reg_0 : DFD1BWP7T port map(CP => clk, D => L1_n_9, Q => L1_col_old_ghost1(0), QN => L1_n_27);
  L1_L3a_L4_row_number_out_reg_2 : EDFKCND1BWP7T port map(CP => clk, CN => L1_n_0, D => L1_n_181, E => L1_n_5, Q => L1_row_old_ghost1(2), QN => L1_n_26);
  L1_L3a_L4_row_number_out_reg_1 : DFD1BWP7T port map(CP => clk, D => L1_n_12, Q => L1_row_old_ghost1(1), QN => L1_n_25);
  L1_L3a_L4_column_number_out_reg_4 : EDFKCND1BWP7T port map(CP => clk, CN => L1_n_0, D => L1_n_184, E => L1_n_1, Q => L1_col_old_ghost1(4), QN => L1_n_20);
  L1_L3a_L4_column_number_out_reg_1 : DFD1BWP7T port map(CP => clk, D => L1_n_10, Q => L1_col_old_ghost1(1), QN => L1_n_19);
  L1_L3a_L4_row_number_out_reg_0 : DFD1BWP7T port map(CP => clk, D => L1_n_11, Q => L1_row_old_ghost1(0), QN => L1_n_18);
  L1_L3a_L4_row_number_out_reg_3 : DFD1BWP7T port map(CP => clk, D => L1_n_13, Q => L1_row_old_ghost1(3), QN => L1_n_16);
  L1_L3a_L4_row_number_out_reg_4 : EDFKCND1BWP7T port map(CP => clk, CN => L1_n_0, D => L1_n_190, E => L1_n_5, Q => L1_row_old_ghost1(4), QN => L1_n_15);
  L1_L1a_g3828 : INVD1BWP7T port map(I => L1_L5_n_14, ZN => L1_L1a_n_180);
  L1_L1a_g9812 : AN4D0BWP7T port map(A1 => L1_L1a_n_179, A2 => L1_L1a_coin_memory(13), A3 => L1_L1a_coin_memory(14), A4 => L1_L1a_coin_memory(15), Z => L1_zero_coins);
  L1_L1a_g9813 : AN4D0BWP7T port map(A1 => L1_L1a_n_178, A2 => L1_L1a_coin_memory(10), A3 => L1_L1a_coin_memory(11), A4 => L1_L1a_coin_memory(12), Z => L1_L1a_n_179);
  L1_L1a_g9814 : AN4D0BWP7T port map(A1 => L1_L1a_n_177, A2 => L1_L1a_coin_memory(6), A3 => L1_L1a_coin_memory(7), A4 => L1_L1a_coin_memory(9), Z => L1_L1a_n_178);
  L1_L1a_g9815 : AN4D0BWP7T port map(A1 => L1_L1a_n_176, A2 => L1_L1a_coin_memory(43), A3 => L1_L1a_coin_memory(4), A4 => L1_L1a_coin_memory(5), Z => L1_L1a_n_177);
  L1_L1a_g9816 : AN4D0BWP7T port map(A1 => L1_L1a_n_175, A2 => L1_L1a_coin_memory(40), A3 => L1_L1a_coin_memory(41), A4 => L1_L1a_coin_memory(42), Z => L1_L1a_n_176);
  L1_L1a_g9817 : AN4D0BWP7T port map(A1 => L1_L1a_n_174, A2 => L1_L1a_coin_memory(37), A3 => L1_L1a_coin_memory(38), A4 => L1_L1a_coin_memory(39), Z => L1_L1a_n_175);
  L1_L1a_g9818 : AN4D0BWP7T port map(A1 => L1_L1a_n_173, A2 => L1_L1a_coin_memory(47), A3 => L1_L1a_coin_memory(8), A4 => L1_L1a_coin_memory(36), Z => L1_L1a_n_174);
  L1_L1a_g9819 : AN4D0BWP7T port map(A1 => L1_L1a_n_172, A2 => L1_L1a_coin_memory(44), A3 => L1_L1a_coin_memory(45), A4 => L1_L1a_coin_memory(46), Z => L1_L1a_n_173);
  L1_L1a_g9820 : CKAN2D1BWP7T port map(A1 => L1_coin_present, A2 => L1_write_coin, Z => score_pulse_int);
  L1_L1a_g9821 : NR3D0BWP7T port map(A1 => L1_L1a_n_171, A2 => L1_L1a_n_162, A3 => L1_L1a_n_134, ZN => L1_coin_present);
  L1_L1a_g9822 : AN4D0BWP7T port map(A1 => L1_L1a_n_169, A2 => L1_L1a_coin_memory(2), A3 => L1_L1a_coin_memory(3), A4 => L1_L1a_coin_memory(35), Z => L1_L1a_n_172);
  L1_L1a_g9823 : OAI221D0BWP7T port map(A1 => L1_L1a_n_147, A2 => L1_L1a_n_206, B1 => L1_L1a_n_195, B2 => L1_L1a_n_138, C => L1_L1a_n_170, ZN => L1_L1a_n_171);
  L1_L1a_g9824 : AOI21D0BWP7T port map(A1 => L1_L1a_n_168, A2 => L1_L1a_n_153, B => L1_L1a_n_159, ZN => L1_L1a_n_170);
  L1_L1a_g9825 : AN4D0BWP7T port map(A1 => L1_L1a_n_167, A2 => L1_L1a_coin_memory(21), A3 => L1_L1a_coin_memory(0), A4 => L1_L1a_coin_memory(1), Z => L1_L1a_n_169);
  L1_L1a_g9826 : AOI211D1BWP7T port map(A1 => L1_L1a_n_136, A2 => L1_L1a_n_104, B => L1_L1a_n_166, C => L1_L1a_n_129, ZN => L1_L1a_n_168);
  L1_L1a_g9827 : AN4D0BWP7T port map(A1 => L1_L1a_n_164, A2 => L1_L1a_coin_memory(23), A3 => L1_L1a_coin_memory(22), A4 => L1_L1a_coin_memory(20), Z => L1_L1a_n_167);
  L1_L1a_g9828 : OAI221D0BWP7T port map(A1 => L1_L1a_n_142, A2 => L1_L1a_n_196, B1 => L1_L1a_n_197, B2 => L1_L1a_n_135, C => L1_L1a_n_165, ZN => L1_L1a_n_166);
  L1_L1a_g9829 : OA221D0BWP7T port map(A1 => L1_L1a_n_113, A2 => L1_L1a_n_203, B1 => L1_L1a_n_183, B2 => L1_L1a_n_202, C => L1_L1a_n_163, Z => L1_L1a_n_165);
  L1_L1a_g9830 : AN4D0BWP7T port map(A1 => L1_L1a_n_161, A2 => L1_L1a_coin_memory(18), A3 => L1_L1a_coin_memory(17), A4 => L1_L1a_coin_memory(16), Z => L1_L1a_n_164);
  L1_L1a_g9831 : AN4D0BWP7T port map(A1 => L1_L1a_n_160, A2 => L1_L1a_n_154, A3 => L1_L1a_n_133, A4 => L1_L1a_n_128, Z => L1_L1a_n_163);
  L1_L1a_g9832 : ND4D0BWP7T port map(A1 => L1_L1a_n_157, A2 => L1_L1a_n_155, A3 => L1_L1a_n_156, A4 => L1_L1a_n_158, ZN => L1_L1a_n_162);
  L1_L1a_g9833 : AN4D0BWP7T port map(A1 => L1_L1a_n_151, A2 => L1_L1a_coin_memory(31), A3 => L1_L1a_coin_memory(19), A4 => L1_L1a_coin_memory(24), Z => L1_L1a_n_161);
  L1_L1a_g9834 : AN4D0BWP7T port map(A1 => L1_L1a_n_152, A2 => L1_L1a_n_150, A3 => L1_L1a_n_139, A4 => L1_L1a_n_115, Z => L1_L1a_n_160);
  L1_L1a_g9835 : OAI221D0BWP7T port map(A1 => L1_L1a_n_145, A2 => L1_L1a_n_194, B1 => L1_L1a_n_193, B2 => L1_L1a_n_119, C => L1_L1a_n_141, ZN => L1_L1a_n_159);
  L1_L1a_g9836 : OA221D0BWP7T port map(A1 => L1_L1a_n_149, A2 => L1_L1a_n_203, B1 => L1_L1a_n_202, B2 => L1_L1a_n_126, C => L1_L1a_n_132, Z => L1_L1a_n_158);
  L1_L1a_g9837 : OA221D0BWP7T port map(A1 => L1_L1a_n_146, A2 => L1_L1a_n_197, B1 => L1_L1a_n_196, B2 => L1_L1a_n_127, C => L1_L1a_n_131, Z => L1_L1a_n_157);
  L1_L1a_g9838 : OA221D0BWP7T port map(A1 => L1_L1a_n_148, A2 => L1_L1a_n_199, B1 => L1_L1a_n_198, B2 => L1_L1a_n_137, C => L1_L1a_n_130, Z => L1_L1a_n_156);
  L1_L1a_g9839 : OA221D0BWP7T port map(A1 => L1_L1a_n_144, A2 => L1_L1a_n_201, B1 => L1_L1a_n_200, B2 => L1_L1a_n_125, C => L1_L1a_n_112, Z => L1_L1a_n_155);
  L1_L1a_g9840 : IAO21D0BWP7T port map(A1 => L1_L1a_n_142, A2 => L1_L1a_n_199, B => L1_L1a_n_140, ZN => L1_L1a_n_154);
  L1_L1a_g9841 : OA22D0BWP7T port map(A1 => L1_L1a_n_143, A2 => L1_L1a_n_200, B1 => L1_L1a_n_201, B2 => L1_L1a_n_116, Z => L1_L1a_n_153);
  L1_L1a_g9842 : OA22D0BWP7T port map(A1 => L1_L1a_n_143, A2 => L1_L1a_n_206, B1 => L1_L1a_n_185, B2 => L1_L1a_n_195, Z => L1_L1a_n_152);
  L1_L1a_g9843 : AN4D0BWP7T port map(A1 => L1_L1a_n_109, A2 => L1_L1a_coin_memory(28), A3 => L1_L1a_coin_memory(29), A4 => L1_L1a_coin_memory(30), Z => L1_L1a_n_151);
  L1_L1a_g9844 : OAI21D0BWP7T port map(A1 => L1_L1a_n_136, A2 => L1_L1a_n_93, B => L1_L1a_n_106, ZN => L1_L1a_n_150);
  L1_L1a_g9845 : CKAN2D1BWP7T port map(A1 => L1_L1a_n_123, A2 => L1_L1a_n_124, Z => L1_L1a_n_149);
  L1_L1a_g9846 : CKAN2D1BWP7T port map(A1 => L1_L1a_n_110, A2 => L1_L1a_n_122, Z => L1_L1a_n_148);
  L1_L1a_g9847 : CKAN2D1BWP7T port map(A1 => L1_L1a_n_111, A2 => L1_L1a_n_121, Z => L1_L1a_n_147);
  L1_L1a_g9848 : CKAN2D1BWP7T port map(A1 => L1_L1a_n_120, A2 => L1_L1a_n_107, Z => L1_L1a_n_146);
  L1_L1a_g9849 : CKAN2D1BWP7T port map(A1 => L1_L1a_n_108, A2 => L1_L1a_n_118, Z => L1_L1a_n_145);
  L1_L1a_g9850 : AOI221D0BWP7T port map(A1 => L1_L1a_n_99, A2 => L1_L1a_coin_memory(41), B1 => L1_L1a_n_91, B2 => L1_L1a_coin_memory(40), C => L1_L1a_n_117, ZN => L1_L1a_n_144);
  L1_L1a_g9851 : AOI32D1BWP7T port map(A1 => L1_L1a_n_105, A2 => L1_L1a_n_84, A3 => L1_L1a_coin_memory(7), B1 => L1_L1a_n_114, B2 => L1_L1a_coin_memory(14), ZN => L1_L1a_n_141);
  L1_L1a_g9852 : AOI21D0BWP7T port map(A1 => L1_L1a_n_198, A2 => L1_L1a_n_195, B => L1_L1a_n_135, ZN => L1_L1a_n_140);
  L1_L1a_g9853 : AO21D0BWP7T port map(A1 => L1_L1a_n_181, A2 => L1_L1a_n_113, B => L1_L1a_n_193, Z => L1_L1a_n_139);
  L1_L1a_g9854 : AOI222D0BWP7T port map(A1 => L1_L1a_n_100, A2 => L1_L1a_coin_memory(6), B1 => L1_L1a_n_99, B2 => L1_L1a_coin_memory(5), C1 => L1_L1a_n_91, C2 => L1_L1a_coin_memory(4), ZN => L1_L1a_n_138);
  L1_L1a_g9855 : AOI222D0BWP7T port map(A1 => L1_L1a_n_100, A2 => L1_L1a_coin_memory(22), B1 => L1_L1a_n_99, B2 => L1_L1a_coin_memory(21), C1 => L1_L1a_n_91, C2 => L1_L1a_coin_memory(20), ZN => L1_L1a_n_137);
  L1_L1a_g9856 : AN3D1BWP7T port map(A1 => L1_L1a_n_113, A2 => L1_L1a_n_187, A3 => L1_L1a_n_204, Z => L1_L1a_n_143);
  L1_L1a_g9857 : AN3D1BWP7T port map(A1 => L1_L1a_n_113, A2 => L1_L1a_n_189, A3 => L1_L1a_n_185, Z => L1_L1a_n_142);
  L1_L1a_g9858 : INR3D0BWP7T port map(A1 => L1_L1a_coin_memory(47), B1 => L1_L1a_n_204, B2 => L1_L1a_n_200, ZN => L1_L1a_n_134);
  L1_L1a_g9859 : AO21D0BWP7T port map(A1 => L1_L1a_n_188, A2 => L1_L1a_n_185, B => L1_L1a_n_201, Z => L1_L1a_n_133);
  L1_L1a_g9860 : IND3D1BWP7T port map(A1 => L1_L1a_n_196, B1 => L1_L1a_coin_memory(31), B2 => L1_L1a_n_84, ZN => L1_L1a_n_132);
  L1_L1a_g9861 : IND3D0BWP7T port map(A1 => L1_L1a_n_198, B1 => L1_L1a_coin_memory(23), B2 => L1_L1a_n_84, ZN => L1_L1a_n_131);
  L1_L1a_g9862 : IND3D1BWP7T port map(A1 => L1_L1a_n_193, B1 => L1_L1a_coin_memory(15), B2 => L1_L1a_n_98, ZN => L1_L1a_n_130);
  L1_L1a_g9863 : AOI21D0BWP7T port map(A1 => L1_L1a_n_181, A2 => L1_L1a_n_192, B => L1_L1a_n_203, ZN => L1_L1a_n_129);
  L1_L1a_g9864 : AO21D0BWP7T port map(A1 => L1_L1a_n_198, A2 => L1_L1a_n_197, B => L1_L1a_n_185, Z => L1_L1a_n_128);
  L1_L1a_g9865 : AOI222D0BWP7T port map(A1 => L1_L1a_n_98, A2 => L1_L1a_coin_memory(30), B1 => L1_L1a_n_91, B2 => L1_L1a_coin_memory(28), C1 => L1_L1a_n_92, C2 => L1_L1a_coin_memory(29), ZN => L1_L1a_n_127);
  L1_L1a_g9866 : ND3D0BWP7T port map(A1 => L1_L1a_n_191, A2 => L1_L1a_n_182, A3 => L1_L1a_n_190, ZN => L1_L1a_n_136);
  L1_L1a_g9867 : CKAN2D1BWP7T port map(A1 => L1_L1a_n_116, A2 => L1_L1a_n_188, Z => L1_L1a_n_135);
  L1_L1a_g9868 : AOI222D0BWP7T port map(A1 => L1_L1a_n_102, A2 => L1_L1a_coin_memory(38), B1 => L1_L1a_n_94, B2 => L1_L1a_coin_memory(36), C1 => L1_L1a_n_93, C2 => L1_L1a_coin_memory(37), ZN => L1_L1a_n_126);
  L1_L1a_g9869 : AOI222D0BWP7T port map(A1 => L1_L1a_n_98, A2 => L1_L1a_coin_memory(46), B1 => L1_L1a_n_86, B2 => L1_L1a_coin_memory(44), C1 => L1_L1a_n_92, C2 => L1_L1a_coin_memory(45), ZN => L1_L1a_n_125);
  L1_L1a_g9870 : AOI22D0BWP7T port map(A1 => L1_L1a_n_92, A2 => L1_L1a_coin_memory(32), B1 => L1_L1a_n_103, B2 => L1_L1a_coin_memory(34), ZN => L1_L1a_n_124);
  L1_L1a_g9871 : AOI22D0BWP7T port map(A1 => L1_L1a_n_101, A2 => L1_L1a_coin_memory(33), B1 => L1_L1a_n_98, B2 => L1_L1a_coin_memory(35), ZN => L1_L1a_n_123);
  L1_L1a_g9872 : AOI22D0BWP7T port map(A1 => L1_L1a_n_98, A2 => L1_L1a_coin_memory(18), B1 => L1_L1a_n_92, B2 => L1_L1a_coin_memory(17), ZN => L1_L1a_n_122);
  L1_L1a_g9873 : AOI22D0BWP7T port map(A1 => L1_L1a_n_98, A2 => L1_L1a_coin_memory(2), B1 => L1_L1a_n_95, B2 => L1_L1a_coin_memory(3), ZN => L1_L1a_n_121);
  L1_L1a_g9874 : AOI22D0BWP7T port map(A1 => L1_L1a_n_99, A2 => L1_L1a_coin_memory(25), B1 => L1_L1a_n_100, B2 => L1_L1a_coin_memory(26), ZN => L1_L1a_n_120);
  L1_L1a_g9875 : AOI22D0BWP7T port map(A1 => L1_L1a_n_101, A2 => L1_L1a_coin_memory(13), B1 => L1_L1a_n_92, B2 => L1_L1a_coin_memory(12), ZN => L1_L1a_n_119);
  L1_L1a_g9876 : AOI22D0BWP7T port map(A1 => L1_L1a_n_102, A2 => L1_L1a_coin_memory(10), B1 => L1_L1a_n_93, B2 => L1_L1a_coin_memory(9), ZN => L1_L1a_n_118);
  L1_L1a_g9877 : AO22D0BWP7T port map(A1 => L1_L1a_n_84, A2 => L1_L1a_coin_memory(43), B1 => L1_L1a_coin_memory(42), B2 => L1_L1a_n_100, Z => L1_L1a_n_117);
  L1_L1a_g9878 : CKND1BWP7T port map(I => L1_L1a_n_114, ZN => L1_L1a_n_115);
  L1_L1a_g9879 : IND3D1BWP7T port map(A1 => L1_L1a_n_182, B1 => L1_L1a_coin_memory(39), B2 => L1_L1a_n_104, ZN => L1_L1a_n_112);
  L1_L1a_g9880 : NR2XD0BWP7T port map(A1 => L1_L1a_n_100, A2 => L1_L1a_n_84, ZN => L1_L1a_n_116);
  L1_L1a_g9881 : NR2D1BWP7T port map(A1 => L1_L1a_n_192, A2 => L1_L1a_n_193, ZN => L1_L1a_n_114);
  L1_L1a_g9882 : NR2XD0BWP7T port map(A1 => L1_L1a_n_98, A2 => L1_L1a_n_92, ZN => L1_L1a_n_113);
  L1_L1a_g9883 : AOI22D0BWP7T port map(A1 => L1_L1a_n_86, A2 => L1_L1a_coin_memory(0), B1 => L1_L1a_n_92, B2 => L1_L1a_coin_memory(1), ZN => L1_L1a_n_111);
  L1_L1a_g9884 : AOI22D0BWP7T port map(A1 => L1_L1a_n_91, A2 => L1_L1a_coin_memory(16), B1 => L1_L1a_n_84, B2 => L1_L1a_coin_memory(19), ZN => L1_L1a_n_110);
  L1_L1a_g9885 : AN4D0BWP7T port map(A1 => L1_L1a_n_75, A2 => L1_L1a_coin_memory(25), A3 => L1_L1a_coin_memory(26), A4 => L1_L1a_coin_memory(27), Z => L1_L1a_n_109);
  L1_L1a_g9886 : AOI22D0BWP7T port map(A1 => L1_L1a_n_94, A2 => L1_L1a_coin_memory(8), B1 => L1_L1a_n_85, B2 => L1_L1a_coin_memory(11), ZN => L1_L1a_n_108);
  L1_L1a_g9887 : AOI22D0BWP7T port map(A1 => L1_L1a_n_91, A2 => L1_L1a_coin_memory(24), B1 => L1_L1a_n_84, B2 => L1_L1a_coin_memory(27), ZN => L1_L1a_n_107);
  L1_L1a_g9888 : INVD0BWP7T port map(I => L1_L1a_n_106, ZN => L1_L1a_n_194);
  L1_L1a_g9889 : INVD0BWP7T port map(I => L1_L1a_n_195, ZN => L1_L1a_n_105);
  L1_L1a_g9890 : INVD0BWP7T port map(I => L1_L1a_n_202, ZN => L1_L1a_n_104);
  L1_L1a_g9891 : NR2D1BWP7T port map(A1 => L1_L1a_n_90, A2 => L1_row_coin(1), ZN => L1_L1a_n_106);
  L1_L1a_g9892 : OR2D1BWP7T port map(A1 => L1_L1a_n_97, A2 => L1_row_coin(1), Z => L1_L1a_n_199);
  L1_L1a_g9893 : OR2D1BWP7T port map(A1 => L1_L1a_n_89, A2 => L1_row_coin(1), Z => L1_L1a_n_201);
  L1_L1a_g9894 : ND2D1BWP7T port map(A1 => L1_L1a_n_88, A2 => L1_L1a_n_65, ZN => L1_L1a_n_203);
  L1_L1a_g9895 : IND2D1BWP7T port map(A1 => L1_L1a_n_89, B1 => L1_row_coin(1), ZN => L1_L1a_n_200);
  L1_L1a_g9896 : ND2D1BWP7T port map(A1 => L1_L1a_n_96, A2 => L1_row_coin(1), ZN => L1_L1a_n_195);
  L1_L1a_g9898 : ND2D1BWP7T port map(A1 => L1_L1a_n_88, A2 => L1_row_coin(1), ZN => L1_L1a_n_202);
  L1_L1a_g9899 : IND2D1BWP7T port map(A1 => L1_L1a_n_97, B1 => L1_row_coin(1), ZN => L1_L1a_n_198);
  L1_L1a_g9900 : INVD1BWP7T port map(I => L1_L1a_n_103, ZN => L1_L1a_n_192);
  L1_L1a_g9901 : INVD0BWP7T port map(I => L1_L1a_n_191, ZN => L1_L1a_n_102);
  L1_L1a_g9902 : INVD0BWP7T port map(I => L1_L1a_n_101, ZN => L1_L1a_n_181);
  L1_L1a_g9903 : INVD1BWP7T port map(I => L1_L1a_n_184, ZN => L1_L1a_n_100);
  L1_L1a_g9904 : INVD0BWP7T port map(I => L1_L1a_n_99, ZN => L1_L1a_n_188);
  L1_L1a_g9905 : INVD1BWP7T port map(I => L1_L1a_n_186, ZN => L1_L1a_n_98);
  L1_L1a_g9906 : ND2D1BWP7T port map(A1 => L1_L1a_n_96, A2 => L1_L1a_n_65, ZN => L1_L1a_n_206);
  L1_L1a_g9907 : ND2D1BWP7T port map(A1 => L1_L1a_n_87, A2 => L1_row_coin(1), ZN => L1_L1a_n_196);
  L1_L1a_g9908 : ND2D1BWP7T port map(A1 => L1_L1a_n_87, A2 => L1_L1a_n_65, ZN => L1_L1a_n_197);
  L1_L1a_g9909 : NR3D0BWP7T port map(A1 => L1_L1a_n_79, A2 => L1_L1a_n_66, A3 => L1_col_coin(0), ZN => L1_L1a_n_103);
  L1_L1a_g9910 : IND3D1BWP7T port map(A1 => L1_col_coin(2), B1 => L1_col_coin(4), B2 => L1_L1a_n_82, ZN => L1_L1a_n_191);
  L1_L1a_g9911 : NR3D0BWP7T port map(A1 => L1_L1a_n_83, A2 => L1_col_coin(1), A3 => L1_L1a_n_67, ZN => L1_L1a_n_101);
  L1_L1a_g9912 : IND3D1BWP7T port map(A1 => L1_L1a_n_79, B1 => L1_col_coin(0), B2 => L1_col_coin(1), ZN => L1_L1a_n_184);
  L1_L1a_g9913 : NR3D0BWP7T port map(A1 => L1_L1a_n_83, A2 => L1_col_coin(1), A3 => L1_col_coin(0), ZN => L1_L1a_n_99);
  L1_L1a_g9914 : IND3D1BWP7T port map(A1 => L1_col_coin(2), B1 => L1_col_coin(4), B2 => L1_L1a_n_80, ZN => L1_L1a_n_186);
  L1_L1a_g9915 : INVD0BWP7T port map(I => L1_L1a_n_204, ZN => L1_L1a_n_95);
  L1_L1a_g9916 : INVD0BWP7T port map(I => L1_L1a_n_190, ZN => L1_L1a_n_94);
  L1_L1a_g9917 : INVD1BWP7T port map(I => L1_L1a_n_183, ZN => L1_L1a_n_93);
  L1_L1a_g9919 : INVD1BWP7T port map(I => L1_L1a_n_185, ZN => L1_L1a_n_91);
  L1_L1a_g9920 : ND2D1BWP7T port map(A1 => L1_L1a_n_78, A2 => L1_row_coin(3), ZN => L1_L1a_n_97);
  L1_L1a_g9921 : INR2D1BWP7T port map(A1 => L1_L1a_n_78, B1 => L1_row_coin(3), ZN => L1_L1a_n_96);
  L1_L1a_g9922 : IND2D1BWP7T port map(A1 => L1_L1a_n_72, B1 => L1_L1a_n_82, ZN => L1_L1a_n_204);
  L1_L1a_g9923 : IND2D1BWP7T port map(A1 => L1_L1a_n_81, B1 => L1_L1a_n_68, ZN => L1_L1a_n_190);
  L1_L1a_g9924 : ND2D1BWP7T port map(A1 => L1_L1a_n_80, A2 => L1_L1a_n_70, ZN => L1_L1a_n_183);
  L1_L1a_g9925 : NR2D1BWP7T port map(A1 => L1_L1a_n_69, A2 => L1_L1a_n_81, ZN => L1_L1a_n_92);
  L1_L1a_g9926 : CKND2D1BWP7T port map(A1 => L1_L1a_n_68, A2 => L1_L1a_n_80, ZN => L1_L1a_n_185);
  L1_L1a_g9928 : INVD0BWP7T port map(I => L1_L1a_n_187, ZN => L1_L1a_n_86);
  L1_L1a_g9929 : INVD0BWP7T port map(I => L1_L1a_n_182, ZN => L1_L1a_n_85);
  L1_L1a_g9930 : CKND1BWP7T port map(I => L1_L1a_n_84, ZN => L1_L1a_n_189);
  L1_L1a_g9931 : IND3D1BWP7T port map(A1 => L1_row_coin(3), B1 => L1_row_coin(2), B2 => L1_L1a_n_71, ZN => L1_L1a_n_90);
  L1_L1a_g9932 : ND2D1BWP7T port map(A1 => L1_L1a_n_76, A2 => L1_row_coin(2), ZN => L1_L1a_n_89);
  L1_L1a_g9933 : NR2XD0BWP7T port map(A1 => L1_L1a_n_77, A2 => L1_row_coin(2), ZN => L1_L1a_n_88);
  L1_L1a_g9934 : IINR4D0BWP7T port map(A1 => L1_row_coin(3), A2 => L1_row_coin(2), B1 => L1_row_coin(4), B2 => L1_row_coin(0), ZN => L1_L1a_n_87);
  L1_L1a_g9935 : ND3D0BWP7T port map(A1 => L1_L1a_n_68, A2 => L1_L1a_n_74, A3 => L1_col_coin(1), ZN => L1_L1a_n_187);
  L1_L1a_g9936 : IND2D1BWP7T port map(A1 => L1_L1a_n_72, B1 => L1_L1a_n_80, ZN => L1_L1a_n_182);
  L1_L1a_g9937 : NR2XD0BWP7T port map(A1 => L1_L1a_n_72, A2 => L1_L1a_n_81, ZN => L1_L1a_n_84);
  L1_L1a_g9938 : ND2D1BWP7T port map(A1 => L1_L1a_n_68, A2 => L1_col_coin(3), ZN => L1_L1a_n_83);
  L1_L1a_g9939 : AN2D1BWP7T port map(A1 => L1_L1a_n_73, A2 => L1_L1a_n_66, Z => L1_L1a_n_82);
  L1_L1a_g9940 : ND2D1BWP7T port map(A1 => L1_L1a_n_73, A2 => L1_col_coin(1), ZN => L1_L1a_n_81);
  L1_L1a_g9941 : AN2D1BWP7T port map(A1 => L1_L1a_n_74, A2 => L1_L1a_n_66, Z => L1_L1a_n_80);
  L1_L1a_g9942 : INVD0BWP7T port map(I => L1_L1a_n_76, ZN => L1_L1a_n_77);
  L1_L1a_g9943 : AN3D0BWP7T port map(A1 => L1_L1a_coin_memory(33), A2 => L1_L1a_coin_memory(32), A3 => L1_L1a_coin_memory(34), Z => L1_L1a_n_75);
  L1_L1a_g9944 : ND2D1BWP7T port map(A1 => L1_L1a_n_70, A2 => L1_col_coin(3), ZN => L1_L1a_n_79);
  L1_L1a_g9945 : INR2XD0BWP7T port map(A1 => L1_L1a_n_71, B1 => L1_row_coin(2), ZN => L1_L1a_n_78);
  L1_L1a_g9946 : INR3D0BWP7T port map(A1 => L1_row_coin(4), B1 => L1_row_coin(0), B2 => L1_row_coin(3), ZN => L1_L1a_n_76);
  L1_L1a_g9947 : NR2D1BWP7T port map(A1 => L1_col_coin(3), A2 => L1_L1a_n_67, ZN => L1_L1a_n_74);
  L1_L1a_g9948 : NR2XD0BWP7T port map(A1 => L1_col_coin(3), A2 => L1_col_coin(0), ZN => L1_L1a_n_73);
  L1_L1a_g9949 : ND2D1BWP7T port map(A1 => L1_col_coin(4), A2 => L1_col_coin(2), ZN => L1_L1a_n_72);
  L1_L1a_g9950 : INVD1BWP7T port map(I => L1_L1a_n_70, ZN => L1_L1a_n_69);
  L1_L1a_g9951 : INR2XD0BWP7T port map(A1 => L1_row_coin(0), B1 => L1_row_coin(4), ZN => L1_L1a_n_71);
  L1_L1a_g9952 : INR2XD0BWP7T port map(A1 => L1_col_coin(2), B1 => L1_col_coin(4), ZN => L1_L1a_n_70);
  L1_L1a_g9953 : NR2XD0BWP7T port map(A1 => L1_col_coin(4), A2 => L1_col_coin(2), ZN => L1_L1a_n_68);
  L1_L1a_g9954 : INVD0BWP7T port map(I => L1_col_coin(0), ZN => L1_L1a_n_67);
  L1_L1a_g9955 : INVD1BWP7T port map(I => L1_col_coin(1), ZN => L1_L1a_n_66);
  L1_L1a_g9957 : INVD1BWP7T port map(I => L1_row_coin(1), ZN => L1_L1a_n_65);
  L1_L1a_g2 : IND2D1BWP7T port map(A1 => L1_L1a_n_90, B1 => L1_row_coin(1), ZN => L1_L1a_n_193);
  L1_L1a_coin_memory_reg_0 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_18, Q => L1_L1a_coin_memory(0));
  L1_L1a_coin_memory_reg_1 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_48, Q => L1_L1a_coin_memory(1));
  L1_L1a_coin_memory_reg_2 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_46, Q => L1_L1a_coin_memory(2));
  L1_L1a_coin_memory_reg_3 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_19, Q => L1_L1a_coin_memory(3));
  L1_L1a_coin_memory_reg_4 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_36, Q => L1_L1a_coin_memory(4));
  L1_L1a_coin_memory_reg_5 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_39, Q => L1_L1a_coin_memory(5));
  L1_L1a_coin_memory_reg_6 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_34, Q => L1_L1a_coin_memory(6));
  L1_L1a_coin_memory_reg_7 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_33, Q => L1_L1a_coin_memory(7));
  L1_L1a_coin_memory_reg_8 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_28, Q => L1_L1a_coin_memory(8));
  L1_L1a_coin_memory_reg_9 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_27, Q => L1_L1a_coin_memory(9));
  L1_L1a_coin_memory_reg_10 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_63, Q => L1_L1a_coin_memory(10));
  L1_L1a_coin_memory_reg_11 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_61, Q => L1_L1a_coin_memory(11));
  L1_L1a_coin_memory_reg_12 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_59, Q => L1_L1a_coin_memory(12));
  L1_L1a_coin_memory_reg_13 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_24, Q => L1_L1a_coin_memory(13));
  L1_L1a_coin_memory_reg_14 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_21, Q => L1_L1a_coin_memory(14));
  L1_L1a_coin_memory_reg_15 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_56, Q => L1_L1a_coin_memory(15));
  L1_L1a_coin_memory_reg_16 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_55, Q => L1_L1a_coin_memory(16));
  L1_L1a_coin_memory_reg_17 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_54, Q => L1_L1a_coin_memory(17));
  L1_L1a_coin_memory_reg_18 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_53, Q => L1_L1a_coin_memory(18));
  L1_L1a_coin_memory_reg_19 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_52, Q => L1_L1a_coin_memory(19));
  L1_L1a_coin_memory_reg_20 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_51, Q => L1_L1a_coin_memory(20));
  L1_L1a_coin_memory_reg_21 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_50, Q => L1_L1a_coin_memory(21));
  L1_L1a_coin_memory_reg_22 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_64, Q => L1_L1a_coin_memory(22));
  L1_L1a_coin_memory_reg_23 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_47, Q => L1_L1a_coin_memory(23));
  L1_L1a_coin_memory_reg_24 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_45, Q => L1_L1a_coin_memory(24));
  L1_L1a_coin_memory_reg_25 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_44, Q => L1_L1a_coin_memory(25));
  L1_L1a_coin_memory_reg_26 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_43, Q => L1_L1a_coin_memory(26));
  L1_L1a_coin_memory_reg_27 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_42, Q => L1_L1a_coin_memory(27));
  L1_L1a_coin_memory_reg_28 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_41, Q => L1_L1a_coin_memory(28));
  L1_L1a_coin_memory_reg_29 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_40, Q => L1_L1a_coin_memory(29));
  L1_L1a_coin_memory_reg_30 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_38, Q => L1_L1a_coin_memory(30));
  L1_L1a_coin_memory_reg_31 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_37, Q => L1_L1a_coin_memory(31));
  L1_L1a_coin_memory_reg_32 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_35, Q => L1_L1a_coin_memory(32));
  L1_L1a_coin_memory_reg_33 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_20, Q => L1_L1a_coin_memory(33));
  L1_L1a_coin_memory_reg_34 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_17, Q => L1_L1a_coin_memory(34));
  L1_L1a_coin_memory_reg_35 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_32, Q => L1_L1a_coin_memory(35));
  L1_L1a_coin_memory_reg_36 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_31, Q => L1_L1a_coin_memory(36));
  L1_L1a_coin_memory_reg_37 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_30, Q => L1_L1a_coin_memory(37));
  L1_L1a_coin_memory_reg_38 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_29, Q => L1_L1a_coin_memory(38));
  L1_L1a_coin_memory_reg_39 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_26, Q => L1_L1a_coin_memory(39));
  L1_L1a_coin_memory_reg_40 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_25, Q => L1_L1a_coin_memory(40));
  L1_L1a_coin_memory_reg_41 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_49, Q => L1_L1a_coin_memory(41));
  L1_L1a_coin_memory_reg_42 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_62, Q => L1_L1a_coin_memory(42));
  L1_L1a_coin_memory_reg_43 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_60, Q => L1_L1a_coin_memory(43));
  L1_L1a_coin_memory_reg_44 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_22, Q => L1_L1a_coin_memory(44));
  L1_L1a_coin_memory_reg_45 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_58, Q => L1_L1a_coin_memory(45));
  L1_L1a_coin_memory_reg_46 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_57, Q => L1_L1a_coin_memory(46));
  L1_L1a_coin_memory_reg_47 : DFQD1BWP7T port map(CP => clk, D => L1_L1a_n_23, Q => L1_L1a_coin_memory(47));
  L1_L1a_g4886 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_11, A2 => L1_L1a_n_198, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(22), ZN => L1_L1a_n_64);
  L1_L1a_g4887 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_9, A2 => L1_L1a_n_191, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(10), ZN => L1_L1a_n_63);
  L1_L1a_g4888 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_11, A2 => L1_L1a_n_201, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(42), ZN => L1_L1a_n_62);
  L1_L1a_g4889 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_9, A2 => L1_L1a_n_182, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(11), ZN => L1_L1a_n_61);
  L1_L1a_g4890 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_14, A2 => L1_L1a_n_201, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(43), ZN => L1_L1a_n_60);
  L1_L1a_g4891 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_224, A2 => L1_L1a_n_193, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(12), ZN => L1_L1a_n_59);
  L1_L1a_g4892 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_224, A2 => L1_L1a_n_200, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(45), ZN => L1_L1a_n_58);
  L1_L1a_g4893 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_16, A2 => L1_L1a_n_200, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(46), ZN => L1_L1a_n_57);
  L1_L1a_g4894 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_16, A2 => L1_L1a_n_193, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(15), ZN => L1_L1a_n_56);
  L1_L1a_g4895 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_13, A2 => L1_L1a_n_199, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(16), ZN => L1_L1a_n_55);
  L1_L1a_g4896 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_224, A2 => L1_L1a_n_199, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(17), ZN => L1_L1a_n_54);
  L1_L1a_g4897 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_16, A2 => L1_L1a_n_199, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(18), ZN => L1_L1a_n_53);
  L1_L1a_g4898 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_14, A2 => L1_L1a_n_199, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(19), ZN => L1_L1a_n_52);
  L1_L1a_g4899 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_13, A2 => L1_L1a_n_198, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(20), ZN => L1_L1a_n_51);
  L1_L1a_g4900 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_10, A2 => L1_L1a_n_198, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(21), ZN => L1_L1a_n_50);
  L1_L1a_g4901 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_10, A2 => L1_L1a_n_201, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(41), ZN => L1_L1a_n_49);
  L1_L1a_g4910 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_224, A2 => L1_L1a_n_206, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(1), ZN => L1_L1a_n_48);
  L1_L1a_g4911 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_14, A2 => L1_L1a_n_198, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(23), ZN => L1_L1a_n_47);
  L1_L1a_g4912 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_16, A2 => L1_L1a_n_206, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(2), ZN => L1_L1a_n_46);
  L1_L1a_g4913 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_13, A2 => L1_L1a_n_197, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(24), ZN => L1_L1a_n_45);
  L1_L1a_g4914 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_10, A2 => L1_L1a_n_197, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(25), ZN => L1_L1a_n_44);
  L1_L1a_g4915 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_11, A2 => L1_L1a_n_197, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(26), ZN => L1_L1a_n_43);
  L1_L1a_g4916 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_14, A2 => L1_L1a_n_197, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(27), ZN => L1_L1a_n_42);
  L1_L1a_g4917 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_13, A2 => L1_L1a_n_196, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(28), ZN => L1_L1a_n_41);
  L1_L1a_g4918 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_224, A2 => L1_L1a_n_196, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(29), ZN => L1_L1a_n_40);
  L1_L1a_g4919 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_10, A2 => L1_L1a_n_195, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(5), ZN => L1_L1a_n_39);
  L1_L1a_g4920 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_16, A2 => L1_L1a_n_196, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(30), ZN => L1_L1a_n_38);
  L1_L1a_g4921 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_14, A2 => L1_L1a_n_196, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(31), ZN => L1_L1a_n_37);
  L1_L1a_g4922 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_13, A2 => L1_L1a_n_195, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(4), ZN => L1_L1a_n_36);
  L1_L1a_g4923 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_224, A2 => L1_L1a_n_203, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(32), ZN => L1_L1a_n_35);
  L1_L1a_g4924 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_11, A2 => L1_L1a_n_195, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(6), ZN => L1_L1a_n_34);
  L1_L1a_g4925 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_14, A2 => L1_L1a_n_195, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(7), ZN => L1_L1a_n_33);
  L1_L1a_g4926 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_16, A2 => L1_L1a_n_203, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(35), ZN => L1_L1a_n_32);
  L1_L1a_g4927 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_12, A2 => L1_L1a_n_190, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(36), ZN => L1_L1a_n_31);
  L1_L1a_g4928 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_12, A2 => L1_L1a_n_183, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(37), ZN => L1_L1a_n_30);
  L1_L1a_g4929 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_12, A2 => L1_L1a_n_191, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(38), ZN => L1_L1a_n_29);
  L1_L1a_g4930 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_9, A2 => L1_L1a_n_190, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(8), ZN => L1_L1a_n_28);
  L1_L1a_g4931 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_9, A2 => L1_L1a_n_183, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(9), ZN => L1_L1a_n_27);
  L1_L1a_g4932 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_12, A2 => L1_L1a_n_182, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(39), ZN => L1_L1a_n_26);
  L1_L1a_g4933 : MOAI22D0BWP7T port map(A1 => L1_L1a_n_13, A2 => L1_L1a_n_201, B1 => L1_L1a_n_180, B2 => L1_L1a_coin_memory(40), ZN => L1_L1a_n_25);
  L1_L1a_g4934 : OAI31D0BWP7T port map(A1 => L1_L1a_n_181, A2 => L1_L1a_n_193, A3 => L1_L1a_n_225, B => L1_L1a_n_6, ZN => L1_L1a_n_24);
  L1_L1a_g4935 : OAI31D0BWP7T port map(A1 => L1_L1a_n_204, A2 => L1_L1a_n_200, A3 => L1_L1a_n_225, B => L1_L1a_n_7, ZN => L1_L1a_n_23);
  L1_L1a_g4936 : OAI31D0BWP7T port map(A1 => L1_L1a_n_187, A2 => L1_L1a_n_200, A3 => L1_L1a_n_225, B => L1_L1a_n_1, ZN => L1_L1a_n_22);
  L1_L1a_g4937 : OAI31D0BWP7T port map(A1 => L1_L1a_n_192, A2 => L1_L1a_n_193, A3 => L1_L1a_n_225, B => L1_L1a_n_8, ZN => L1_L1a_n_21);
  L1_L1a_g4938 : OAI31D0BWP7T port map(A1 => L1_L1a_n_181, A2 => L1_L1a_n_203, A3 => L1_L1a_n_225, B => L1_L1a_n_3, ZN => L1_L1a_n_20);
  L1_L1a_g4939 : OAI31D0BWP7T port map(A1 => L1_L1a_n_204, A2 => L1_L1a_n_206, A3 => L1_L1a_n_225, B => L1_L1a_n_0, ZN => L1_L1a_n_19);
  L1_L1a_g4940 : OAI31D0BWP7T port map(A1 => L1_L1a_n_187, A2 => L1_L1a_n_206, A3 => L1_L1a_n_225, B => L1_L1a_n_2, ZN => L1_L1a_n_18);
  L1_L1a_g4941 : OAI31D0BWP7T port map(A1 => L1_L1a_n_192, A2 => L1_L1a_n_203, A3 => L1_L1a_n_225, B => L1_L1a_n_5, ZN => L1_L1a_n_17);
  L1_L1a_g4942 : OR2D1BWP7T port map(A1 => L1_L1a_n_225, A2 => L1_L1a_n_186, Z => L1_L1a_n_16);
  L1_L1a_g4944 : OR2D1BWP7T port map(A1 => L1_L1a_n_225, A2 => L1_L1a_n_189, Z => L1_L1a_n_14);
  L1_L1a_g4945 : OR2D1BWP7T port map(A1 => L1_L1a_n_225, A2 => L1_L1a_n_185, Z => L1_L1a_n_13);
  L1_L1a_g4946 : OR2D1BWP7T port map(A1 => L1_L1a_n_225, A2 => L1_L1a_n_202, Z => L1_L1a_n_12);
  L1_L1a_g4947 : OR2D1BWP7T port map(A1 => L1_L1a_n_225, A2 => L1_L1a_n_184, Z => L1_L1a_n_11);
  L1_L1a_g4948 : OR2D1BWP7T port map(A1 => L1_L1a_n_225, A2 => L1_L1a_n_188, Z => L1_L1a_n_10);
  L1_L1a_g4949 : OR2D1BWP7T port map(A1 => L1_L1a_n_225, A2 => L1_L1a_n_194, Z => L1_L1a_n_9);
  L1_L1a_g4950 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(14), ZN => L1_L1a_n_8);
  L1_L1a_g4951 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(47), ZN => L1_L1a_n_7);
  L1_L1a_g4952 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(13), ZN => L1_L1a_n_6);
  L1_L1a_g4953 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(34), ZN => L1_L1a_n_5);
  L1_L1a_g4954 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(33), ZN => L1_L1a_n_3);
  L1_L1a_g4955 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(0), ZN => L1_L1a_n_2);
  L1_L1a_g4956 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(44), ZN => L1_L1a_n_1);
  L1_L1a_g4957 : ND2D1BWP7T port map(A1 => L1_L1a_n_180, A2 => L1_L1a_coin_memory(3), ZN => L1_L1a_n_0);
  L1_L1a_g9958 : IND2D1BWP7T port map(A1 => L1_L1a_n_225, B1 => L1_L1a_n_92, ZN => L1_L1a_n_224);
  L1_L1a_g9959 : ND2D1BWP7T port map(A1 => L1_write_coin, A2 => L1_L1a_n_180, ZN => L1_L1a_n_225);
  L1_L1b_g182 : AO22D0BWP7T port map(A1 => L1_col_new_pacman(3), A2 => L1_L1b_n_0, B1 => L1_n_23, B2 => xcoordinates_int(3), Z => L1_col_coin(3));
  L1_L1b_g183 : AO22D0BWP7T port map(A1 => L1_L1b_n_0, A2 => L1_row_new_pacman(1), B1 => L1_n_23, B2 => ycoordinates_int(1), Z => L1_row_coin(1));
  L1_L1b_g184 : AO22D0BWP7T port map(A1 => L1_row_new_pacman(4), A2 => L1_L1b_n_0, B1 => L1_n_23, B2 => ycoordinates_int(4), Z => L1_row_coin(4));
  L1_L1b_g185 : AO22D0BWP7T port map(A1 => L1_L1b_n_0, A2 => L1_col_new_pacman(2), B1 => L1_n_23, B2 => xcoordinates_int(2), Z => L1_col_coin(2));
  L1_L1b_g186 : AO22D0BWP7T port map(A1 => L1_L1b_n_0, A2 => L1_row_new_pacman(0), B1 => L1_n_23, B2 => ycoordinates_int(0), Z => L1_row_coin(0));
  L1_L1b_g187 : AO22D0BWP7T port map(A1 => L1_row_new_pacman(3), A2 => L1_L1b_n_0, B1 => L1_n_23, B2 => ycoordinates_int(3), Z => L1_row_coin(3));
  L1_L1b_g188 : AO22D0BWP7T port map(A1 => L1_L1b_n_0, A2 => L1_col_new_pacman(0), B1 => L1_n_23, B2 => xcoordinates_int(0), Z => L1_col_coin(0));
  L1_L1b_g189 : AO22D0BWP7T port map(A1 => L1_L1b_n_0, A2 => L1_col_new_pacman(1), B1 => L1_n_23, B2 => xcoordinates_int(1), Z => L1_col_coin(1));
  L1_L1b_g190 : AO22D0BWP7T port map(A1 => L1_L1b_n_0, A2 => L1_row_new_pacman(2), B1 => L1_n_23, B2 => ycoordinates_int(2), Z => L1_row_coin(2));
  L1_L1b_g191 : AO22D0BWP7T port map(A1 => L1_col_new_pacman(4), A2 => L1_L1b_n_0, B1 => L1_n_23, B2 => xcoordinates_int(4), Z => L1_col_coin(4));
  L1_L1b_g192 : INVD1BWP7T port map(I => L1_n_23, ZN => L1_L1b_n_0);
  L1_L3b_g256 : NR2D1BWP7T port map(A1 => L1_L3b_n_5, A2 => L1_L3b_n_6, ZN => L1_ghost2_map_select);
  L1_L3b_g307 : AO21D0BWP7T port map(A1 => L1_pos_is_wall, A2 => L1_L3b_n_0, B => L1_L3b_n_1, Z => L1_L3b_n_2);
  L1_L3b_L5_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => L1_L3b_n_0, Q => L1_L3b_n_6);
  L1_L3b_g309 : INR4D0BWP7T port map(A1 => L1_ghost2_start, B1 => L1_L3b_n_6, B2 => L1_L3b_L5_state(0), B3 => game_over_out_int, ZN => L1_L3b_n_1);
  L1_L3b_g310 : NR3D0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3b_n_5, A3 => L1_L3b_n_6, ZN => L1_L3b_n_0);
  L1_L3b_L5_state_reg_0 : DFD1BWP7T port map(CP => clk, D => L1_L3b_n_2, Q => L1_L3b_L5_state(0), QN => L1_L3b_n_5);
  L1_L3c_g1491 : OAI222D0BWP7T port map(A1 => L1_L3c_n_59, A2 => L1_L3c_n_46, B1 => L1_L3c_n_43, B2 => L1_L3c_n_60, C1 => L1_L3c_n_44, C2 => L1_L3c_n_16, ZN => L1_row_new_pacman(4));
  L1_L3c_g1492 : OAI222D0BWP7T port map(A1 => L1_L3c_n_59, A2 => L1_L3c_n_32, B1 => L1_L3c_n_34, B2 => L1_L3c_n_60, C1 => L1_L3c_n_40, C2 => L1_L3c_n_15, ZN => L1_col_new_pacman(4));
  L1_L3c_g1493 : OAI21D0BWP7T port map(A1 => L1_L3c_n_55, A2 => L1_L3c_n_34, B => L1_L3c_n_61, ZN => L1_col_new_pacman(3));
  L1_L3c_g1494 : OAI222D0BWP7T port map(A1 => L1_L3c_n_58, A2 => L1_L3c_n_46, B1 => L1_L3c_n_43, B2 => L1_L3c_n_55, C1 => L1_L3c_n_44, C2 => L1_L3c_n_14, ZN => L1_row_new_pacman(3));
  L1_L3c_g1495 : MAOI22D0BWP7T port map(A1 => L1_col_old_pacman(3), A2 => L1_L3c_n_41, B1 => L1_L3c_n_58, B2 => L1_L3c_n_32, ZN => L1_L3c_n_61);
  L1_L3c_g1496 : MAOI22D0BWP7T port map(A1 => L1_L3c_n_53, A2 => L1_L3c_n_25, B1 => L1_L3c_n_53, B2 => L1_L3c_n_25, ZN => L1_L3c_n_60);
  L1_L3c_g1497 : MAOI22D0BWP7T port map(A1 => L1_L3c_n_57, A2 => L1_L3c_n_30, B1 => L1_L3c_n_57, B2 => L1_L3c_n_30, ZN => L1_L3c_n_59);
  L1_L3c_g1498 : HA1D0BWP7T port map(A => L1_L3c_n_26, B => L1_L3c_n_49, CO => L1_L3c_n_57, S => L1_L3c_n_58);
  L1_L3c_g1499 : OAI21D0BWP7T port map(A1 => L1_L3c_n_51, A2 => L1_L3c_n_43, B => L1_L3c_n_54, ZN => L1_row_new_pacman(2));
  L1_L3c_g1500 : OAI21D0BWP7T port map(A1 => L1_L3c_n_51, A2 => L1_L3c_n_34, B => L1_L3c_n_56, ZN => L1_col_new_pacman(2));
  L1_L3c_g1501 : AOI22D0BWP7T port map(A1 => L1_L3c_n_52, A2 => L1_L3c_n_31, B1 => L1_col_old_pacman(2), B2 => L1_L3c_n_41, ZN => L1_L3c_n_56);
  L1_L3c_g1502 : AOI22D0BWP7T port map(A1 => L1_L3c_n_52, A2 => L1_L3c_n_47, B1 => L1_row_old_pacman(2), B2 => L1_L3c_n_45, ZN => L1_L3c_n_54);
  L1_L3c_g1503 : MAOI22D0BWP7T port map(A1 => L1_L3c_n_48, A2 => L1_L3c_n_24, B1 => L1_L3c_n_48, B2 => L1_L3c_n_24, ZN => L1_L3c_n_55);
  L1_L3c_g1504 : INR2XD0BWP7T port map(A1 => L1_L3c_n_48, B1 => L1_L3c_n_24, ZN => L1_L3c_n_53);
  L1_L3c_g1505 : OAI21D0BWP7T port map(A1 => L1_L3c_n_38, A2 => L1_L3c_n_34, B => L1_L3c_n_50, ZN => L1_col_new_pacman(1));
  L1_L3c_g1506 : OAI222D0BWP7T port map(A1 => L1_L3c_n_39, A2 => L1_L3c_n_46, B1 => L1_L3c_n_43, B2 => L1_L3c_n_38, C1 => L1_L3c_n_44, C2 => L1_L3c_n_18, ZN => L1_row_new_pacman(1));
  L1_L3c_g1507 : AO222D0BWP7T port map(A1 => L1_L3c_n_42, A2 => L1_L3c_n_21, B1 => L1_L3c_n_47, B2 => L1_L3c_n_27, C1 => L1_row_old_pacman(0), C2 => L1_L3c_n_45, Z => L1_row_new_pacman(0));
  L1_L3c_g1508 : AO222D0BWP7T port map(A1 => L1_L3c_n_33, A2 => L1_L3c_n_21, B1 => L1_L3c_n_31, B2 => L1_L3c_n_27, C1 => L1_col_old_pacman(0), C2 => L1_L3c_n_41, Z => L1_col_new_pacman(0));
  L1_L3c_g1509 : AO21D0BWP7T port map(A1 => L1_L3c_n_36, A2 => L1_L3c_n_29, B => L1_L3c_n_49, Z => L1_L3c_n_52);
  L1_L3c_g1510 : MAOI22D0BWP7T port map(A1 => L1_col_old_pacman(1), A2 => L1_L3c_n_41, B1 => L1_L3c_n_39, B2 => L1_L3c_n_32, ZN => L1_L3c_n_50);
  L1_L3c_g1511 : MAOI22D0BWP7T port map(A1 => L1_L3c_n_35, A2 => L1_L3c_n_22, B1 => L1_L3c_n_35, B2 => L1_L3c_n_22, ZN => L1_L3c_n_51);
  L1_L3c_g1512 : NR2XD0BWP7T port map(A1 => L1_L3c_n_36, A2 => L1_L3c_n_29, ZN => L1_L3c_n_49);
  L1_L3c_g1513 : INR2XD0BWP7T port map(A1 => L1_L3c_n_35, B1 => L1_L3c_n_22, ZN => L1_L3c_n_48);
  L1_L3c_g1514 : CKND1BWP7T port map(I => L1_L3c_n_46, ZN => L1_L3c_n_47);
  L1_L3c_g1515 : IND3D0BWP7T port map(A1 => L1_L3c_move(3), B1 => L1_L3c_move(1), B2 => L1_L3c_n_37, ZN => L1_L3c_n_46);
  L1_L3c_g1516 : CKND1BWP7T port map(I => L1_L3c_n_44, ZN => L1_L3c_n_45);
  L1_L3c_g1517 : CKND1BWP7T port map(I => L1_L3c_n_43, ZN => L1_L3c_n_42);
  L1_L3c_g1518 : AOI211D0BWP7T port map(A1 => L1_L3c_move(3), A2 => L1_L3c_move(1), B => L1_L3c_n_19, C => L1_L3c_n_20, ZN => L1_L3c_n_44);
  L1_L3c_g1519 : IND3D0BWP7T port map(A1 => L1_L3c_move(1), B1 => L1_L3c_move(3), B2 => L1_L3c_n_37, ZN => L1_L3c_n_43);
  L1_L3c_g1520 : CKND1BWP7T port map(I => L1_L3c_n_41, ZN => L1_L3c_n_40);
  L1_L3c_g1521 : OAI211D0BWP7T port map(A1 => L1_L3c_n_17, A2 => L1_L3c_n_13, B => L1_L3c_n_20, C => L1_L3c_n_19, ZN => L1_L3c_n_41);
  L1_L3c_g1522 : OA21D0BWP7T port map(A1 => L1_L3c_n_27, A2 => L1_L3c_n_28, B => L1_L3c_n_36, Z => L1_L3c_n_39);
  L1_L3c_g1523 : XNR2D1BWP7T port map(A1 => L1_L3c_n_21, A2 => L1_L3c_n_23, ZN => L1_L3c_n_38);
  L1_L3c_g1524 : CKND1BWP7T port map(I => L1_L3c_n_20, ZN => L1_L3c_n_37);
  L1_L3c_g1525 : ND2D1BWP7T port map(A1 => L1_L3c_n_28, A2 => L1_L3c_n_27, ZN => L1_L3c_n_36);
  L1_L3c_g1526 : NR2XD0BWP7T port map(A1 => L1_L3c_n_21, A2 => L1_L3c_n_23, ZN => L1_L3c_n_35);
  L1_L3c_g1527 : CKND1BWP7T port map(I => L1_L3c_n_34, ZN => L1_L3c_n_33);
  L1_L3c_g1528 : CKND1BWP7T port map(I => L1_L3c_n_32, ZN => L1_L3c_n_31);
  L1_L3c_g1529 : ND3D0BWP7T port map(A1 => L1_L3c_n_19, A2 => L1_L3c_n_13, A3 => L1_L3c_move(0), ZN => L1_L3c_n_34);
  L1_L3c_g1530 : ND3D0BWP7T port map(A1 => L1_L3c_n_19, A2 => L1_L3c_n_17, A3 => L1_L3c_move(2), ZN => L1_L3c_n_32);
  L1_L3c_g1531 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(3), A2 => L1_L3c_n_13, B1 => L1_col_old_pacman(3), B2 => L1_L3c_move(2), ZN => L1_L3c_n_26);
  L1_L3c_g1532 : OAI22D0BWP7T port map(A1 => L1_row_old_pacman(4), A2 => L1_L3c_move(2), B1 => L1_col_old_pacman(4), B2 => L1_L3c_n_13, ZN => L1_L3c_n_30);
  L1_L3c_g1533 : AO22D0BWP7T port map(A1 => L1_row_old_pacman(2), A2 => L1_L3c_n_13, B1 => L1_L3c_move(2), B2 => L1_col_old_pacman(2), Z => L1_L3c_n_29);
  L1_L3c_g1534 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(1), A2 => L1_L3c_n_13, B1 => L1_col_old_pacman(1), B2 => L1_L3c_move(2), ZN => L1_L3c_n_28);
  L1_L3c_g1535 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(0), A2 => L1_L3c_n_13, B1 => L1_col_old_pacman(0), B2 => L1_L3c_move(2), ZN => L1_L3c_n_27);
  L1_L3c_g1536 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(4), A2 => L1_L3c_move(3), B1 => L1_col_old_pacman(4), B2 => L1_L3c_move(0), ZN => L1_L3c_n_25);
  L1_L3c_g1537 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(3), A2 => L1_L3c_move(3), B1 => L1_col_old_pacman(3), B2 => L1_L3c_move(0), ZN => L1_L3c_n_24);
  L1_L3c_g1538 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(1), A2 => L1_L3c_move(3), B1 => L1_col_old_pacman(1), B2 => L1_L3c_move(0), ZN => L1_L3c_n_23);
  L1_L3c_g1539 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(2), A2 => L1_L3c_move(3), B1 => L1_col_old_pacman(2), B2 => L1_L3c_move(0), ZN => L1_L3c_n_22);
  L1_L3c_g1540 : AOI22D0BWP7T port map(A1 => L1_row_old_pacman(0), A2 => L1_L3c_move(3), B1 => L1_col_old_pacman(0), B2 => L1_L3c_move(0), ZN => L1_L3c_n_21);
  L1_L3c_g1541 : ND2D0BWP7T port map(A1 => L1_L3c_n_13, A2 => L1_L3c_n_17, ZN => L1_L3c_n_20);
  L1_L3c_g1542 : NR2D0BWP7T port map(A1 => L1_L3c_move(3), A2 => L1_L3c_move(1), ZN => L1_L3c_n_19);
  L1_L3c_g1544 : INVD0BWP7T port map(I => L1_L3c_move(0), ZN => L1_L3c_n_17);
  L1_L3c_g1548 : INVD1BWP7T port map(I => L1_L3c_move(2), ZN => L1_L3c_n_13);
  L1_L3c_CR1_column_number_out_reg_2 : DFQD1BWP7T port map(CP => clk, D => L1_L3c_n_5, Q => L1_col_old_pacman(2));
  L1_L3c_CR1_row_number_out_reg_0 : DFQD1BWP7T port map(CP => clk, D => L1_L3c_n_7, Q => L1_row_old_pacman(0));
  L1_L3c_CR1_row_number_out_reg_2 : DFQD1BWP7T port map(CP => clk, D => L1_L3c_n_4, Q => L1_row_old_pacman(2));
  L1_L3c_CR1_column_number_out_reg_1 : DFQD1BWP7T port map(CP => clk, D => L1_L3c_n_8, Q => L1_col_old_pacman(1));
  L1_L3c_CR1_column_number_out_reg_0 : DFQD1BWP7T port map(CP => clk, D => L1_L3c_n_12, Q => L1_col_old_pacman(0));
  L1_L3c_CR1_column_number_out_reg_3 : DFQD1BWP7T port map(CP => clk, D => L1_L3c_n_11, Q => L1_col_old_pacman(3));
  L1_L3c_g475 : AO221D0BWP7T port map(A1 => L1_L3c_n_0, A2 => L1_col_old_pacman(0), B1 => L1_write_coin, B2 => L1_col_new_pacman(0), C => game_over_out_int, Z => L1_L3c_n_12);
  L1_L3c_g476 : AO221D0BWP7T port map(A1 => L1_L3c_n_0, A2 => L1_col_old_pacman(3), B1 => L1_col_new_pacman(3), B2 => L1_write_coin, C => game_over_out_int, Z => L1_L3c_n_11);
  L1_L3c_g477 : AO221D0BWP7T port map(A1 => L1_L3c_n_0, A2 => L1_row_old_pacman(4), B1 => L1_row_new_pacman(4), B2 => L1_write_coin, C => game_over_out_int, Z => L1_L3c_n_10);
  L1_L3c_g478 : AO221D0BWP7T port map(A1 => L1_L3c_n_0, A2 => L1_row_old_pacman(1), B1 => L1_write_coin, B2 => L1_row_new_pacman(1), C => game_over_out_int, Z => L1_L3c_n_9);
  L1_L3c_g479 : AO221D0BWP7T port map(A1 => L1_L3c_n_0, A2 => L1_col_old_pacman(1), B1 => L1_write_coin, B2 => L1_col_new_pacman(1), C => game_over_out_int, Z => L1_L3c_n_8);
  L1_L3c_g480 : AO22D0BWP7T port map(A1 => L1_L3c_n_1, A2 => L1_row_old_pacman(0), B1 => L1_row_new_pacman(0), B2 => L1_L3c_n_2, Z => L1_L3c_n_7);
  L1_L3c_g481 : AO22D0BWP7T port map(A1 => L1_L3c_n_1, A2 => L1_col_old_pacman(4), B1 => L1_col_new_pacman(4), B2 => L1_L3c_n_2, Z => L1_L3c_n_6);
  L1_L3c_g482 : AO22D0BWP7T port map(A1 => L1_L3c_n_1, A2 => L1_col_old_pacman(2), B1 => L1_col_new_pacman(2), B2 => L1_L3c_n_2, Z => L1_L3c_n_5);
  L1_L3c_g483 : AO22D0BWP7T port map(A1 => L1_L3c_n_1, A2 => L1_row_old_pacman(2), B1 => L1_row_new_pacman(2), B2 => L1_L3c_n_2, Z => L1_L3c_n_4);
  L1_L3c_g484 : AO22D0BWP7T port map(A1 => L1_L3c_n_1, A2 => L1_row_old_pacman(3), B1 => L1_row_new_pacman(3), B2 => L1_L3c_n_2, Z => L1_L3c_n_3);
  L1_L3c_g485 : NR2D1BWP7T port map(A1 => game_over_out_int, A2 => L1_L3c_n_0, ZN => L1_L3c_n_2);
  L1_L3c_g486 : NR2XD0BWP7T port map(A1 => game_over_out_int, A2 => L1_write_coin, ZN => L1_L3c_n_1);
  L1_L3c_g487 : INVD1BWP7T port map(I => L1_write_coin, ZN => L1_L3c_n_0);
  L1_L3c_CR1_row_number_out_reg_1 : DFD1BWP7T port map(CP => clk, D => L1_L3c_n_9, Q => L1_row_old_pacman(1), QN => L1_L3c_n_18);
  L1_L3c_CR1_row_number_out_reg_4 : DFD1BWP7T port map(CP => clk, D => L1_L3c_n_10, Q => L1_row_old_pacman(4), QN => L1_L3c_n_16);
  L1_L3c_CR1_column_number_out_reg_4 : DFD1BWP7T port map(CP => clk, D => L1_L3c_n_6, Q => L1_col_old_pacman(4), QN => L1_L3c_n_15);
  L1_L3c_CR1_row_number_out_reg_3 : DFD1BWP7T port map(CP => clk, D => L1_L3c_n_3, Q => L1_row_old_pacman(3), QN => L1_L3c_n_14);
  L1_L3c_PC1_g171 : ND2D1BWP7T port map(A1 => L1_L3c_PC1_n_8, A2 => L1_L3c_PC1_n_9, ZN => L1_pacman_ready);
  L1_L3c_PC1_g172 : NR2XD0BWP7T port map(A1 => L1_L3c_PC1_n_7, A2 => L1_L3c_PC1_state(1), ZN => L1_pacman_map_select);
  L1_L3c_PC1_g317 : MOAI22D0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3c_PC1_n_2, B1 => L1_pos_is_wall, B2 => L1_L3c_PC1_n_3, ZN => L1_L3c_PC1_n_5);
  L1_L3c_PC1_g318 : NR3D0BWP7T port map(A1 => L1_L3c_PC1_n_1, A2 => game_over_out_int, A3 => L1_L3c_PC1_state(1), ZN => L1_L3c_PC1_n_4);
  L1_L3c_PC1_g319 : INR4D0BWP7T port map(A1 => L1_L3c_PC1_n_9, B1 => L1_L3c_PC1_n_7, B2 => L1_pacman_dead, B3 => game_over_out_int, ZN => L1_L3c_PC1_n_3);
  L1_L3c_PC1_g320 : ND4D0BWP7T port map(A1 => L1_pacman_start, A2 => L1_L3c_PC1_n_9, A3 => L1_L3c_PC1_n_7, A4 => L1_L3c_PC1_n_8, ZN => L1_L3c_PC1_n_2);
  L1_L3c_PC1_g321 : OAI21D0BWP7T port map(A1 => L1_pos_is_wall, A2 => L1_pacman_dead, B => L1_L3c_PC1_state(0), ZN => L1_L3c_PC1_n_1);
  L1_L3c_PC1_g322 : INVD0BWP7T port map(I => L1_pos_is_wall, ZN => L1_L3c_PC1_n_0);
  L1_L3c_PC1_state_reg_0 : DFD1BWP7T port map(CP => clk, D => L1_L3c_PC1_n_5, Q => L1_L3c_PC1_state(0), QN => L1_L3c_PC1_n_7);
  L1_L3c_PC1_state_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => L1_L3c_PC1_n_3, D => L1_L3c_PC1_n_0, Q => L1_write_coin, QN => L1_L3c_PC1_n_8);
  L1_L3c_PC1_state_reg_1 : DFD1BWP7T port map(CP => clk, D => L1_L3c_PC1_n_4, Q => L1_L3c_PC1_state(1), QN => L1_L3c_PC1_n_9);
  L1_L2_g2 : OR2D1BWP7T port map(A1 => L1_L2_c_g1, A2 => L1_L2_c_g2, Z => L1_pacman_dead);
  L1_L2_IB1_g329 : NR4D0BWP7T port map(A1 => L1_L2_IB1_n_11, A2 => L1_L2_IB1_n_4, A3 => L1_L2_IB1_n_9, A4 => L1_L2_IB1_n_0, ZN => L1_L2_c_g1);
  L1_L2_IB1_g330 : ND4D0BWP7T port map(A1 => L1_L2_IB1_n_10, A2 => L1_L2_IB1_n_1, A3 => L1_L2_IB1_n_8, A4 => L1_L2_IB1_n_5, ZN => L1_L2_IB1_n_11);
  L1_L2_IB1_g331 : NR4D0BWP7T port map(A1 => L1_L2_IB1_n_7, A2 => L1_L2_IB1_n_3, A3 => L1_L2_IB1_n_2, A4 => L1_L2_IB1_n_6, ZN => L1_L2_IB1_n_10);
  L1_L2_IB1_g332 : MAOI22D0BWP7T port map(A1 => L1_row_old_pacman(4), A2 => L1_row_old_ghost1(4), B1 => L1_row_old_pacman(4), B2 => L1_row_old_ghost1(4), ZN => L1_L2_IB1_n_9);
  L1_L2_IB1_g333 : XNR2D1BWP7T port map(A1 => L1_col_old_pacman(0), A2 => L1_col_old_ghost1(0), ZN => L1_L2_IB1_n_8);
  L1_L2_IB1_g334 : CKXOR2D0BWP7T port map(A1 => L1_row_old_pacman(0), A2 => L1_row_old_ghost1(0), Z => L1_L2_IB1_n_7);
  L1_L2_IB1_g335 : CKXOR2D0BWP7T port map(A1 => L1_col_old_pacman(1), A2 => L1_col_old_ghost1(1), Z => L1_L2_IB1_n_6);
  L1_L2_IB1_g336 : MOAI22D0BWP7T port map(A1 => L1_row_old_pacman(1), A2 => L1_row_old_ghost1(1), B1 => L1_row_old_pacman(1), B2 => L1_row_old_ghost1(1), ZN => L1_L2_IB1_n_5);
  L1_L2_IB1_g337 : MAOI22D0BWP7T port map(A1 => L1_row_old_pacman(2), A2 => L1_row_old_ghost1(2), B1 => L1_row_old_pacman(2), B2 => L1_row_old_ghost1(2), ZN => L1_L2_IB1_n_4);
  L1_L2_IB1_g338 : CKXOR2D0BWP7T port map(A1 => L1_col_old_pacman(3), A2 => L1_col_old_ghost1(3), Z => L1_L2_IB1_n_3);
  L1_L2_IB1_g339 : CKXOR2D0BWP7T port map(A1 => L1_col_old_pacman(4), A2 => L1_col_old_ghost1(4), Z => L1_L2_IB1_n_2);
  L1_L2_IB1_g340 : XNR2D1BWP7T port map(A1 => L1_col_old_pacman(2), A2 => L1_col_old_ghost1(2), ZN => L1_L2_IB1_n_1);
  L1_L2_IB1_g341 : MAOI22D0BWP7T port map(A1 => L1_row_old_pacman(3), A2 => L1_row_old_ghost1(3), B1 => L1_row_old_pacman(3), B2 => L1_row_old_ghost1(3), ZN => L1_L2_IB1_n_0);
  L1_L2_IB2_g149 : NR4D0BWP7T port map(A1 => L1_L2_IB2_n_0, A2 => L1_L2_IB2_n_1, A3 => L1_row_old_pacman(1), A4 => L1_row_old_pacman(0), ZN => L1_L2_c_g2);
  L1_L2_IB2_g150 : IIND4D0BWP7T port map(A1 => L1_col_old_pacman(0), A2 => L1_row_old_pacman(4), B1 => L1_row_old_pacman(2), B2 => L1_row_old_pacman(3), ZN => L1_L2_IB2_n_1);
  L1_L2_IB2_g151 : IIND4D0BWP7T port map(A1 => L1_col_old_pacman(4), A2 => L1_col_old_pacman(1), B1 => L1_col_old_pacman(2), B2 => L1_col_old_pacman(3), ZN => L1_L2_IB2_n_0);
  L1_L6a_LBL1_g1129 : AO22D0BWP7T port map(A1 => L1_L6a_LBL1_n_57, A2 => L1_L6a_LBL1_state(1), B1 => L1_L6a_LBL1_n_54, B2 => L1_L6a_LBL1_n_62, Z => L1_pacman_start);
  L1_L6a_LBL1_g1130 : OAI22D0BWP7T port map(A1 => L1_L6a_LBL1_n_56, A2 => L1_L6a_LBL1_state(3), B1 => L1_L6a_LBL1_n_65, B2 => L1_L6a_LBL1_state(2), ZN => L1_L6a_c_rst_int);
  L1_L6a_LBL1_g1131 : NR2XD0BWP7T port map(A1 => L1_L6a_LBL1_n_53, A2 => L1_L6a_LBL1_state(2), ZN => L1_ghost1_start);
  L1_L6a_LBL1_g1132 : NR4D0BWP7T port map(A1 => L1_L6a_LBL1_n_55, A2 => L1_L6a_LBL1_state(0), A3 => L1_L6a_LBL1_state(3), A4 => L1_L6a_LBL1_state(1), ZN => L1_ghost2_start);
  L1_L6a_LBL1_g1133 : NR2XD0BWP7T port map(A1 => L1_L6a_LBL1_n_56, A2 => L1_L6a_LBL1_state(3), ZN => L1_L6a_LBL1_n_57);
  L1_L6a_LBL1_g1134 : INR2D1BWP7T port map(A1 => L1_L6a_LBL1_n_63, B1 => L1_L6a_LBL1_state(1), ZN => L1_L6a_LBL1_n_62);
  L1_L6a_LBL1_g1136 : OAI22D0BWP7T port map(A1 => L1_L6a_LBL1_n_55, A2 => L1_L6a_LBL1_state(0), B1 => L1_L6a_LBL1_n_54, B2 => L1_L6a_LBL1_state(2), ZN => L1_L6a_LBL1_n_56);
  L1_L6a_LBL1_g1137 : ND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_54, A2 => L1_L6a_LBL1_state(1), ZN => L1_L6a_LBL1_n_65);
  L1_L6a_LBL1_g1138 : NR2XD0BWP7T port map(A1 => L1_L6a_LBL1_state(2), A2 => L1_L6a_LBL1_state(3), ZN => L1_L6a_LBL1_n_64);
  L1_L6a_LBL1_g1139 : CKAN2D1BWP7T port map(A1 => L1_L6a_LBL1_state(2), A2 => L1_L6a_LBL1_state(3), Z => L1_L6a_LBL1_n_63);
  L1_L6a_LBL1_g2 : MUX2ND0BWP7T port map(I0 => L1_L6a_LBL1_state(3), I1 => L1_L6a_LBL1_state(0), S => L1_L6a_LBL1_state(1), ZN => L1_L6a_LBL1_n_53);
  L1_L6a_LBL1_state_reg_3 : DFQD1BWP7T port map(CP => clk, D => L1_L6a_LBL1_n_50, Q => L1_L6a_LBL1_state(3));
  L1_L6a_LBL1_g2534 : ND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_51, A2 => L1_L6a_LBL1_n_22, ZN => L1_L6a_LBL1_n_52);
  L1_L6a_LBL1_state_reg_1 : DFXQD1BWP7T port map(CP => clk, DA => L1_L6a_LBL1_n_24, DB => L1_L6a_LBL1_n_48, SA => L1_L6a_LBL1_n_74, Q => L1_L6a_LBL1_state(1));
  L1_L6a_LBL1_g2537 : NR4D0BWP7T port map(A1 => L1_L6a_LBL1_n_43, A2 => L1_L6a_LBL1_n_46, A3 => L1_L6a_LBL1_n_41, A4 => L1_L6a_LBL1_n_25, ZN => L1_L6a_LBL1_n_51);
  L1_L6a_LBL1_g2538 : OAI32D1BWP7T port map(A1 => L1_L6a_LBL1_n_20, A2 => L1_L6a_LBL1_n_74, A3 => L1_L6a_LBL1_n_47, B1 => L1_L6a_LBL1_n_12, B2 => L1_L6a_LBL1_n_36, ZN => L1_L6a_LBL1_n_50);
  L1_L6a_LBL1_g2539 : ND3D0BWP7T port map(A1 => L1_L6a_LBL1_n_45, A2 => L1_L6a_LBL1_n_30, A3 => L1_L6a_LBL1_n_17, ZN => L1_L6a_LBL1_n_49);
  L1_L6a_LBL1_g2540 : INR4D0BWP7T port map(A1 => L1_L6a_LBL1_n_30, B1 => L1_L6a_LBL1_n_25, B2 => L1_L6a_LBL1_n_40, B3 => L1_L6a_LBL1_n_41, ZN => L1_L6a_LBL1_n_48);
  L1_L6a_LBL1_g2541 : OAI211D1BWP7T port map(A1 => L1_L6a_LBL1_n_4, A2 => L1_L6a_LBL1_n_38, B => L1_L6a_LBL1_n_44, C => L1_L6a_LBL1_n_27, ZN => L1_L6a_LBL1_n_47);
  L1_L6a_LBL1_g2542 : OAI21D0BWP7T port map(A1 => L1_L6a_LBL1_n_76, A2 => reset, B => L1_L6a_LBL1_n_42, ZN => L1_L6a_LBL1_n_46);
  L1_L6a_LBL1_g2543 : AOI211XD0BWP7T port map(A1 => L1_L6a_LBL1_n_74, A2 => L1_L6a_LBL1_n_29, B => L1_L6a_LBL1_n_34, C => L1_L6a_LBL1_n_26, ZN => L1_L6a_LBL1_n_45);
  L1_L6a_LBL1_g2544 : CKND1BWP7T port map(I => L1_L6a_LBL1_n_43, ZN => L1_L6a_LBL1_n_44);
  L1_L6a_LBL1_g2545 : ND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_39, A2 => L1_L6a_LBL1_n_35, ZN => L1_L6a_LBL1_n_43);
  L1_L6a_LBL1_g2546 : AOI22D0BWP7T port map(A1 => L1_L6a_LBL1_n_74, A2 => L1_L6a_LBL1_n_15, B1 => L1_L6a_LBL1_n_20, B2 => L1_L6a_LBL1_n_5, ZN => L1_L6a_LBL1_n_42);
  L1_L6a_LBL1_g2547 : NR3D0BWP7T port map(A1 => L1_L6a_LBL1_n_32, A2 => L1_L6a_LBL1_n_9, A3 => L1_L6a_hundredandtwenty, ZN => L1_L6a_LBL1_n_41);
  L1_L6a_LBL1_g2548 : IAO21D0BWP7T port map(A1 => L1_L6a_LBL1_n_33, A2 => reset, B => L1_L6a_LBL1_n_16, ZN => L1_L6a_LBL1_n_40);
  L1_L6a_LBL1_g2549 : AOI33D1BWP7T port map(A1 => L1_L6a_LBL1_n_31, A2 => L1_L6a_LBL1_n_9, A3 => L1_L6a_LBL1_n_4, B1 => L1_L6a_LBL1_n_23, B2 => L1_L6a_hundredandtwenty, B3 => L1_L6a_LBL1_n_4, ZN => L1_L6a_LBL1_n_39);
  L1_L6a_LBL1_g2550 : AOI31D0BWP7T port map(A1 => L1_L6a_eighty, A2 => L1_L6a_LBL1_n_21, A3 => L1_L6a_LBL1_n_2, B => reset, ZN => L1_L6a_LBL1_n_38);
  L1_L6a_LBL1_g2551 : INVD0BWP7T port map(I => L1_L6a_LBL1_n_74, ZN => L1_L6a_LBL1_n_36);
  L1_L6a_LBL1_g2553 : IND4D0BWP7T port map(A1 => reset, B1 => L1_ghost1_ready, B2 => L1_pacman_ready, B3 => L1_L6a_LBL1_n_14, ZN => L1_L6a_LBL1_n_35);
  L1_L6a_LBL1_g2554 : IOA21D1BWP7T port map(A1 => L1_L6a_LBL1_n_20, A2 => L1_pacman_ready, B => L1_L6a_LBL1_n_18, ZN => L1_L6a_LBL1_n_34);
  L1_L6a_LBL1_g2555 : OA22D0BWP7T port map(A1 => L1_L6a_LBL1_n_14, A2 => L1_L6a_LBL1_n_20, B1 => L1_L6a_LBL1_n_3, B2 => L1_L6a_LBL1_n_23, Z => L1_L6a_LBL1_n_33);
  L1_L6a_LBL1_g2556 : ND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_31, A2 => L1_L6a_LBL1_n_4, ZN => L1_L6a_LBL1_n_32);
  L1_L6a_LBL1_g2557 : INR2D1BWP7T port map(A1 => L1_L6a_LBL1_n_23, B1 => L1_L6a_sixty, ZN => L1_L6a_LBL1_n_31);
  L1_L6a_LBL1_g2558 : IND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_63, B1 => L1_L6a_LBL1_n_24, ZN => L1_L6a_LBL1_n_29);
  L1_L6a_LBL1_g2559 : ND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_19, A2 => L1_L6a_LBL1_n_20, ZN => L1_L6a_LBL1_n_30);
  L1_L6a_LBL1_g2561 : IND3D1BWP7T port map(A1 => L1_L6a_LBL1_n_76, B1 => L1_L6a_LBL1_n_16, B2 => L1_L6a_sixty, ZN => L1_L6a_LBL1_n_27);
  L1_L6a_LBL1_g2562 : AOI21D0BWP7T port map(A1 => L1_L6a_eighty, A2 => L1_L6a_LBL1_n_6, B => L1_L6a_LBL1_n_22, ZN => L1_L6a_LBL1_n_26);
  L1_L6a_LBL1_g2563 : NR2D1BWP7T port map(A1 => L1_L6a_LBL1_n_17, A2 => L1_L6a_LBL1_n_5, ZN => L1_L6a_LBL1_n_25);
  L1_L6a_LBL1_g2564 : CKAN2D1BWP7T port map(A1 => L1_L6a_LBL1_n_15, A2 => L1_L6a_LBL1_n_65, Z => L1_L6a_LBL1_n_24);
  L1_L6a_LBL1_g2565 : AN2D1BWP7T port map(A1 => L1_L6a_LBL1_n_14, A2 => L1_L6a_LBL1_n_2, Z => L1_L6a_LBL1_n_23);
  L1_L6a_LBL1_g2566 : INVD1BWP7T port map(I => L1_L6a_LBL1_n_22, ZN => L1_L6a_LBL1_n_21);
  L1_L6a_LBL1_g2567 : AOI211XD0BWP7T port map(A1 => L1_L6a_sixty, A2 => L1_L6a_LBL1_n_3, B => L1_L6a_LBL1_n_6, C => L1_L6a_LBL1_n_5, ZN => L1_L6a_LBL1_n_19);
  L1_L6a_LBL1_g2568 : OAI211D1BWP7T port map(A1 => L1_ghost1_ready, A2 => L1_L6a_hundredandtwenty, B => L1_L6a_LBL1_n_14, C => L1_L6a_LBL1_n_4, ZN => L1_L6a_LBL1_n_18);
  L1_L6a_LBL1_g2569 : ND3D0BWP7T port map(A1 => L1_L6a_LBL1_n_63, A2 => L1_L6a_LBL1_n_8, A3 => L1_L6a_LBL1_state(1), ZN => L1_L6a_LBL1_n_22);
  L1_L6a_LBL1_g2570 : INR3D0BWP7T port map(A1 => L1_L6a_LBL1_n_64, B1 => L1_L6a_LBL1_state(1), B2 => L1_L6a_LBL1_n_7, ZN => L1_L6a_LBL1_n_20);
  L1_L6a_LBL1_g2571 : ND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_62, A2 => L1_L6a_LBL1_n_8, ZN => L1_L6a_LBL1_n_17);
  L1_L6a_LBL1_g2572 : AN2D1BWP7T port map(A1 => L1_L6a_LBL1_n_4, A2 => L1_L6a_LBL1_n_2, Z => L1_L6a_LBL1_n_16);
  L1_L6a_LBL1_g2573 : IAO21D0BWP7T port map(A1 => L1_L6a_LBL1_state(3), A2 => L1_L6a_LBL1_state(0), B => L1_L6a_LBL1_n_64, ZN => L1_L6a_LBL1_n_15);
  L1_L6a_LBL1_g2574 : INR3D0BWP7T port map(A1 => L1_L6a_LBL1_state(2), B1 => L1_L6a_LBL1_state(3), B2 => L1_L6a_LBL1_n_65, ZN => L1_L6a_LBL1_n_14);
  L1_L6a_LBL1_g2575 : AOI21D0BWP7T port map(A1 => L1_L6a_LBL1_state(3), A2 => L1_L6a_LBL1_state(1), B => L1_L6a_LBL1_n_63, ZN => L1_L6a_LBL1_n_12);
  L1_L6a_LBL1_g2576 : OAI21D0BWP7T port map(A1 => L1_L6a_LBL1_state(1), A2 => L1_L6a_LBL1_state(0), B => L1_L6a_LBL1_n_63, ZN => L1_L6a_LBL1_n_11);
  L1_L6a_LBL1_g2577 : IND3D1BWP7T port map(A1 => L1_L6a_LBL1_state(1), B1 => L1_L6a_LBL1_state(0), B2 => L1_L6a_LBL1_n_64, ZN => L1_L6a_LBL1_n_10);
  L1_L6a_LBL1_g2579 : INVD0BWP7T port map(I => L1_L6a_LBL1_n_7, ZN => L1_L6a_LBL1_n_8);
  L1_L6a_LBL1_g2580 : NR2D1BWP7T port map(A1 => L1_L6a_forty, A2 => L1_L6a_eighty, ZN => L1_L6a_LBL1_n_9);
  L1_L6a_LBL1_g2581 : IND2D1BWP7T port map(A1 => reset, B1 => L1_L6a_LBL1_state(0), ZN => L1_L6a_LBL1_n_7);
  L1_L6a_LBL1_g2582 : NR2D1BWP7T port map(A1 => L1_L6a_LBL1_n_3, A2 => L1_ghost1_ready, ZN => L1_L6a_LBL1_n_6);
  L1_L6a_LBL1_g2583 : NR2XD0BWP7T port map(A1 => L1_pacman_ready, A2 => L1_L6a_LBL1_n_2, ZN => L1_L6a_LBL1_n_5);
  L1_L6a_LBL1_g2584 : NR2XD0BWP7T port map(A1 => L1_pacman_ready, A2 => reset, ZN => L1_L6a_LBL1_n_4);
  L1_L6a_LBL1_g2585 : INVD1BWP7T port map(I => L1_pacman_ready, ZN => L1_L6a_LBL1_n_3);
  L1_L6a_LBL1_g2586 : INVD1BWP7T port map(I => L1_ghost1_ready, ZN => L1_L6a_LBL1_n_2);
  L1_L6a_LBL1_g2600 : NR3D0BWP7T port map(A1 => L1_L6a_LBL1_n_14, A2 => L1_L6a_LBL1_n_75, A3 => reset, ZN => L1_L6a_LBL1_n_74);
  L1_L6a_LBL1_g2601 : ND2D1BWP7T port map(A1 => L1_L6a_LBL1_n_10, A2 => L1_L6a_LBL1_n_11, ZN => L1_L6a_LBL1_n_75);
  L1_L6a_LBL1_g2602 : IND2D1BWP7T port map(A1 => L1_L6a_LBL1_state(0), B1 => L1_L6a_LBL1_n_63, ZN => L1_L6a_LBL1_n_76);
  L1_L6a_LBL1_state_reg_2 : DFD1BWP7T port map(CP => clk, D => L1_L6a_LBL1_n_52, Q => L1_L6a_LBL1_state(2), QN => L1_L6a_LBL1_n_55);
  L1_L6a_LBL1_state_reg_0 : DFD1BWP7T port map(CP => clk, D => L1_L6a_LBL1_n_49, Q => L1_L6a_LBL1_state(0), QN => L1_L6a_LBL1_n_54);
  L1_L6a_LBL2_g291 : IND2D1BWP7T port map(A1 => L1_L6a_LBL2_count(5), B1 => L1_L6a_LBL2_n_23, ZN => L1_L6a_forty);
  L1_L6a_LBL2_g292 : IIND4D0BWP7T port map(A1 => L1_L6a_LBL2_n_24, A2 => L1_L6a_LBL2_count(6), B1 => L1_L6a_LBL2_n_22, B2 => L1_L6a_LBL2_n_18, ZN => L1_L6a_sixty);
  L1_L6a_LBL2_g293 : OAI21D0BWP7T port map(A1 => L1_L6a_LBL2_n_20, A2 => L1_L6a_LBL2_n_18, B => L1_L6a_LBL2_n_15, ZN => L1_L6a_hundredandtwenty);
  L1_L6a_LBL2_g294 : IND3D1BWP7T port map(A1 => L1_L6a_LBL2_n_24, B1 => L1_L6a_LBL2_n_15, B2 => L1_L6a_LBL2_n_19, ZN => L1_L6a_eighty);
  L1_L6a_LBL2_g295 : AOI211XD0BWP7T port map(A1 => L1_L6a_LBL2_count(3), A2 => L1_L6a_LBL2_count(4), B => L1_L6a_LBL2_n_21, C => L1_L6a_LBL2_count(6), ZN => L1_L6a_LBL2_n_23);
  L1_L6a_LBL2_g296 : OAI21D0BWP7T port map(A1 => L1_L6a_LBL2_n_16, A2 => L1_L6a_LBL2_count(2), B => L1_L6a_LBL2_count(5), ZN => L1_L6a_LBL2_n_22);
  L1_L6a_LBL2_g297 : INVD1BWP7T port map(I => L1_L6a_LBL2_n_20, ZN => L1_L6a_LBL2_n_21);
  L1_L6a_LBL2_g298 : AO21D0BWP7T port map(A1 => L1_L6a_LBL2_n_17, A2 => L1_L6a_LBL2_n_14, B => L1_L6a_LBL2_n_18, Z => L1_L6a_LBL2_n_19);
  L1_L6a_LBL2_g299 : IND3D1BWP7T port map(A1 => L1_L6a_LBL2_n_17, B1 => L1_L6a_LBL2_count(2), B2 => L1_L6a_LBL2_count(4), ZN => L1_L6a_LBL2_n_20);
  L1_L6a_LBL2_g300 : AN2D1BWP7T port map(A1 => L1_L6a_LBL2_count(5), A2 => L1_L6a_LBL2_count(4), Z => L1_L6a_LBL2_n_24);
  L1_L6a_LBL2_g301 : ND2D1BWP7T port map(A1 => L1_L6a_LBL2_count(5), A2 => L1_L6a_LBL2_count(3), ZN => L1_L6a_LBL2_n_18);
  L1_L6a_LBL2_g302 : AN2D0BWP7T port map(A1 => L1_L6a_LBL2_count(1), A2 => L1_L6a_LBL2_count(0), Z => L1_L6a_LBL2_n_16);
  L1_L6a_LBL2_g304 : NR2XD0BWP7T port map(A1 => L1_L6a_LBL2_count(1), A2 => L1_L6a_LBL2_count(0), ZN => L1_L6a_LBL2_n_17);
  L1_L6a_LBL2_new_count_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L6a_LBL2_n_0, D => L1_L6a_LBL2_n_13, Q => L1_L6a_LBL2_count(5));
  L1_L6a_LBL2_new_count_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L6a_LBL2_n_0, D => L1_L6a_LBL2_n_12, Q => L1_L6a_LBL2_count(3));
  L1_L6a_LBL2_g238 : MOAI22D0BWP7T port map(A1 => L1_L6a_LBL2_n_9, A2 => L1_L6a_LBL2_count(5), B1 => L1_L6a_LBL2_n_9, B2 => L1_L6a_LBL2_count(5), ZN => L1_L6a_LBL2_n_13);
  L1_L6a_LBL2_new_count_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L6a_LBL2_n_0, D => L1_L6a_LBL2_n_10, Q => L1_L6a_LBL2_count(4));
  L1_L6a_LBL2_g241 : MOAI22D0BWP7T port map(A1 => L1_L6a_LBL2_n_6, A2 => L1_L6a_LBL2_count(3), B1 => L1_L6a_LBL2_n_6, B2 => L1_L6a_LBL2_count(3), ZN => L1_L6a_LBL2_n_12);
  L1_L6a_LBL2_g242 : MOAI22D0BWP7T port map(A1 => L1_L6a_LBL2_n_8, A2 => L1_L6a_LBL2_count(6), B1 => L1_L6a_LBL2_n_8, B2 => L1_L6a_LBL2_count(6), ZN => L1_L6a_LBL2_n_11);
  L1_L6a_LBL2_g243 : MOAI22D0BWP7T port map(A1 => L1_L6a_LBL2_n_32, A2 => L1_L6a_LBL2_count(4), B1 => L1_L6a_LBL2_n_32, B2 => L1_L6a_LBL2_count(4), ZN => L1_L6a_LBL2_n_10);
  L1_L6a_LBL2_g244 : IND2D1BWP7T port map(A1 => L1_L6a_LBL2_n_32, B1 => L1_L6a_LBL2_count(4), ZN => L1_L6a_LBL2_n_9);
  L1_L6a_LBL2_new_count_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L6a_LBL2_n_4, D => L1_L6a_LBL2_n_0, Q => L1_L6a_LBL2_count(1));
  L1_L6a_LBL2_g246 : MOAI22D0BWP7T port map(A1 => L1_L6a_LBL2_n_3, A2 => L1_L6a_LBL2_count(2), B1 => L1_L6a_LBL2_n_3, B2 => L1_L6a_LBL2_count(2), ZN => L1_L6a_LBL2_n_7);
  L1_L6a_LBL2_g247 : IND2D1BWP7T port map(A1 => L1_L6a_LBL2_n_32, B1 => L1_L6a_LBL2_n_24, ZN => L1_L6a_LBL2_n_8);
  L1_L6a_LBL2_g248 : IND2D1BWP7T port map(A1 => L1_L6a_LBL2_n_3, B1 => L1_L6a_LBL2_count(2), ZN => L1_L6a_LBL2_n_6);
  L1_L6a_LBL2_new_count_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L6a_LBL2_n_2, D => L1_L6a_LBL2_n_0, Q => L1_L6a_LBL2_count(0));
  L1_L6a_LBL2_g251 : MOAI22D0BWP7T port map(A1 => L1_L6a_LBL2_n_1, A2 => L1_L6a_LBL2_count(1), B1 => L1_L6a_LBL2_n_1, B2 => L1_L6a_LBL2_count(1), ZN => L1_L6a_LBL2_n_4);
  L1_L6a_LBL2_g252 : IND2D1BWP7T port map(A1 => L1_L6a_LBL2_n_1, B1 => L1_L6a_LBL2_count(1), ZN => L1_L6a_LBL2_n_3);
  L1_L6a_LBL2_g253 : CKXOR2D0BWP7T port map(A1 => L1_L6a_LBL2_count(0), A2 => L1_vc_pulse, Z => L1_L6a_LBL2_n_2);
  L1_L6a_LBL2_g254 : ND2D1BWP7T port map(A1 => L1_vc_pulse, A2 => L1_L6a_LBL2_count(0), ZN => L1_L6a_LBL2_n_1);
  L1_L6a_LBL2_g267 : INVD1BWP7T port map(I => L1_L6a_c_rst_int, ZN => L1_L6a_LBL2_n_0);
  L1_L6a_LBL2_new_count_reg_6 : DFKCND1BWP7T port map(CP => clk, CN => L1_L6a_LBL2_n_0, D => L1_L6a_LBL2_n_11, Q => L1_L6a_LBL2_count(6), QN => L1_L6a_LBL2_n_15);
  L1_L6a_LBL2_new_count_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => L1_L6a_LBL2_n_7, D => L1_L6a_LBL2_n_0, Q => L1_L6a_LBL2_count(2), QN => L1_L6a_LBL2_n_14);
  L1_L6a_LBL2_g2 : IND3D1BWP7T port map(A1 => L1_L6a_LBL2_n_3, B1 => L1_L6a_LBL2_count(3), B2 => L1_L6a_LBL2_count(2), ZN => L1_L6a_LBL2_n_32);
  L1_L3a_L0_FF1_data_out_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_ghost1(3), D => L1_L3a_L0_FF1_n_0, Q => L1_L3a_L0_data_intermediate(3));
  L1_L3a_L0_FF1_data_out_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_ghost1(2), D => L1_L3a_L0_FF1_n_0, Q => L1_L3a_L0_data_intermediate(2));
  L1_L3a_L0_FF1_data_out_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_ghost1(0), D => L1_L3a_L0_FF1_n_0, Q => L1_L3a_L0_data_intermediate(0));
  L1_L3a_L0_FF1_data_out_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_ghost1(1), D => L1_L3a_L0_FF1_n_0, Q => L1_L3a_L0_data_intermediate(1));
  L1_L3a_L0_FF1_g7 : INVD1BWP7T port map(I => game_over_out_int, ZN => L1_L3a_L0_FF1_n_0);
  L1_L3a_L0_FF2_data_out_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3a_L0_data_intermediate(3), D => L1_L3a_L0_FF2_n_0, Q => L1_L3a_data_buffed(3));
  L1_L3a_L0_FF2_data_out_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3a_L0_data_intermediate(2), D => L1_L3a_L0_FF2_n_0, Q => L1_L3a_data_buffed(2));
  L1_L3a_L0_FF2_data_out_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3a_L0_data_intermediate(0), D => L1_L3a_L0_FF2_n_0, Q => L1_L3a_data_buffed(0));
  L1_L3a_L0_FF2_data_out_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3a_L0_data_intermediate(1), D => L1_L3a_L0_FF2_n_0, Q => L1_L3a_data_buffed(1));
  L1_L3a_L0_FF2_g7 : INVD1BWP7T port map(I => game_over_out_int, ZN => L1_L3a_L0_FF2_n_0);
  L2_g4918 : AO21D0BWP7T port map(A1 => L2_screencontrol_n_58, A2 => L2_in_st_go_sel, B => reset, Z => L2_score_reset_or);
  L2_g4919 : INR2XD0BWP7T port map(A1 => user_begin, B1 => L2_n_523, ZN => L2_screencontrol_n_58);
  L2_g4920 : IND4D0BWP7T port map(A1 => L2_n_552, B1 => L2_n_515, B2 => L2_n_518, B3 => L2_n_519, ZN => L2_n_523);
  L2_g4921 : IINR4D0BWP7T port map(A1 => L2_n_517, A2 => L2_n_516, B1 => L2_vgacontrol_hcount(1), B2 => L2_vgacontrol_hcount(0), ZN => L2_n_519);
  L2_g4922 : NR4D0BWP7T port map(A1 => L2_vgacontrol_vcount(3), A2 => L2_vgacontrol_vcount(4), A3 => L2_vgacontrol_hcount(9), A4 => L2_vgacontrol_hcount(2), ZN => L2_n_518);
  L2_g4923 : NR4D0BWP7T port map(A1 => L2_vgacontrol_vcount(2), A2 => L2_vgacontrol_vcount(9), A3 => L2_vgacontrol_hcount(4), A4 => L2_vgacontrol_hcount(5), ZN => L2_n_517);
  L2_g4924 : NR4D0BWP7T port map(A1 => L2_vgacontrol_hcount(6), A2 => L2_vgacontrol_hcount(8), A3 => L2_vgacontrol_hcount(7), A4 => L2_vgacontrol_hcount(3), ZN => L2_n_516);
  L2_g4925 : IINR4D0BWP7T port map(A1 => L2_vgacontrol_vcount(7), A2 => L2_vgacontrol_vcount(8), B1 => L2_vgacontrol_vcount(1), B2 => L2_vgacontrol_vcount(0), ZN => L2_n_515);
  L2_g4926 : AN2D1BWP7T port map(A1 => L2_screencontrol_state(0), A2 => L2_screencontrol_state(1), Z => L2_in_st_go_sel);
  L2_g4927 : ND2D1BWP7T port map(A1 => L2_vgacontrol_vcount(5), A2 => L2_vgacontrol_vcount(6), ZN => L2_n_552);
  L2_shift_L12_shift_sync_reg : DFKCNQD1BWP7T port map(CP => clk, CN => L2_calc_start_internal, D => L2_n_283, Q => L2_shift_shift_pulse);
  L2_vgacontrol_in_blue_reg : DFD0BWP7T port map(CP => clk, D => L2_n_507, Q => UNCONNECTED, QN => L2_n_512);
  L2_vgacontrol_in_green_reg : DFD0BWP7T port map(CP => clk, D => L2_n_511, Q => UNCONNECTED0, QN => L2_n_514);
  L2_vgacontrol_in_red_reg : DFD0BWP7T port map(CP => clk, D => L2_n_510, Q => UNCONNECTED1, QN => L2_n_513);
  L2_g12453 : OAI211D1BWP7T port map(A1 => L2_in_go_sprite_type(3), A2 => L2_n_508, B => L2_n_483, C => L2_n_424, ZN => L2_n_541);
  L2_g12455 : INVD4BWP7T port map(I => L2_n_514, ZN => green);
  L2_g12457 : INVD4BWP7T port map(I => L2_n_513, ZN => red);
  L2_g12458 : OR2D1BWP7T port map(A1 => L2_n_509, A2 => L2_n_410, Z => L2_n_545);
  L2_g12459 : IND3D1BWP7T port map(A1 => L2_n_498, B1 => L2_n_415, B2 => L2_n_424, ZN => L2_n_543);
  L2_g12460 : ND4D0BWP7T port map(A1 => L2_n_499, A2 => L2_n_485, A3 => L2_n_424, A4 => L2_n_397, ZN => L2_n_540);
  L2_g12462 : INVD4BWP7T port map(I => L2_n_512, ZN => blue);
  L2_g12463 : AO31D1BWP7T port map(A1 => L2_n_497, A2 => L2_in_go_colour(1), A3 => L2_n_533, B => L2_n_506, Z => L2_n_511);
  L2_g12464 : AO31D1BWP7T port map(A1 => L2_n_497, A2 => L2_in_go_colour(2), A3 => L2_n_533, B => L2_n_505, Z => L2_n_510);
  L2_g12465 : OAI211D1BWP7T port map(A1 => L2_n_271, A2 => L2_n_476, B => L2_n_501, C => L2_n_446, ZN => L2_n_544);
  L2_g12466 : OAI221D0BWP7T port map(A1 => L2_n_416, A2 => L2_n_312, B1 => L2_n_334, B2 => L2_n_291, C => L2_n_503, ZN => L2_n_509);
  L2_g12467 : OAI221D0BWP7T port map(A1 => L2_n_246, A2 => L2_n_292, B1 => L2_n_294, B2 => L2_n_239, C => L2_n_504, ZN => L2_n_550);
  L2_g12468 : AN3D1BWP7T port map(A1 => L2_n_500, A2 => L2_n_533, A3 => L2_vgacontrol_vcount(5), Z => L2_n_537);
  L2_g12469 : OAI222D0BWP7T port map(A1 => L2_n_495, A2 => L2_in_go_sprite_type(4), B1 => L2_n_231, B2 => L2_n_428, C1 => L2_n_250, C2 => L2_n_423, ZN => L2_n_508);
  L2_g12470 : ND4D0BWP7T port map(A1 => L2_n_490, A2 => L2_n_486, A3 => L2_n_424, A4 => L2_n_413, ZN => L2_n_542);
  L2_g12471 : IAO21D0BWP7T port map(A1 => L2_rgb_score(0), A2 => L2_rgb_video(0), B => L2_n_502, ZN => L2_n_507);
  L2_g12472 : IAO21D0BWP7T port map(A1 => L2_rgb_video(1), A2 => L2_rgb_score(2), B => L2_n_502, ZN => L2_n_506);
  L2_g12473 : IAO21D0BWP7T port map(A1 => L2_rgb_video(2), A2 => L2_rgb_score(2), B => L2_n_502, ZN => L2_n_505);
  L2_g12474 : AOI222D0BWP7T port map(A1 => L2_n_492, A2 => L2_score_score_sprite_type(1), B1 => L2_n_456, B2 => L2_n_276, C1 => L2_n_394, C2 => L2_n_267, ZN => L2_n_504);
  L2_g12475 : AOI221D0BWP7T port map(A1 => L2_n_403, A2 => L2_n_263, B1 => L2_n_363, B2 => L2_n_351, C => L2_n_496, ZN => L2_n_503);
  L2_g12476 : AOI211XD0BWP7T port map(A1 => L2_n_303, A2 => L2_n_298, B => L2_n_491, C => L2_n_410, ZN => L2_n_501);
  L2_g12477 : IND4D0BWP7T port map(A1 => L2_n_478, B1 => L2_n_384, B2 => L2_n_471, B3 => L2_n_481, ZN => L2_n_547);
  L2_g12478 : INR4D0BWP7T port map(A1 => L2_n_488, B1 => L2_vgacontrol_vcount(8), B2 => L2_vgacontrol_vcount(9), B3 => L2_n_522, ZN => L2_n_500);
  L2_g12479 : OAI221D0BWP7T port map(A1 => L2_n_300, A2 => L2_n_294, B1 => L2_n_299, B2 => L2_n_229, C => L2_n_494, ZN => L2_n_551);
  L2_g12480 : IND2D1BWP7T port map(A1 => L2_n_533, B1 => L2_n_497, ZN => L2_n_502);
  L2_g12481 : AN4D1BWP7T port map(A1 => L2_n_488, A2 => L2_n_411, A3 => L2_n_356, A4 => L2_vgacontrol_vcount(5), Z => L2_n_535);
  L2_g12482 : IND4D0BWP7T port map(A1 => L2_n_448, B1 => L2_n_471, B2 => L2_n_472, B3 => L2_n_473, ZN => L2_n_548);
  L2_g12483 : IINR4D0BWP7T port map(A1 => L2_n_488, A2 => L2_n_436, B1 => L2_n_533, B2 => L2_vgacontrol_vcount(9), ZN => L2_n_536);
  L2_g12484 : OA21D0BWP7T port map(A1 => L2_n_443, A2 => L2_n_312, B => L2_n_493, Z => L2_n_499);
  L2_g12485 : OAI222D0BWP7T port map(A1 => L2_n_479, A2 => L2_n_272, B1 => L2_n_262, B2 => L2_n_454, C1 => L2_n_271, C2 => L2_n_467, ZN => L2_n_498);
  L2_g12486 : IND3D1BWP7T port map(A1 => L2_n_477, B1 => L2_n_455, B2 => L2_n_475, ZN => L2_n_549);
  L2_g12487 : OAI222D0BWP7T port map(A1 => L2_n_469, A2 => L2_n_272, B1 => L2_n_438, B2 => L2_n_466, C1 => L2_n_297, C2 => L2_n_332, ZN => L2_n_496);
  L2_g12488 : NR3D0BWP7T port map(A1 => L2_n_482, A2 => L2_vgacontrol_vcount(9), A3 => L2_vgacontrol_hcount(9), ZN => L2_n_497);
  L2_g12489 : AOI221D0BWP7T port map(A1 => L2_n_360, A2 => L2_n_308, B1 => L2_n_289, B2 => L2_n_284, C => L2_n_489, ZN => L2_n_495);
  L2_g12490 : AOI31D0BWP7T port map(A1 => L2_n_464, A2 => L2_n_439, A3 => L2_score_score_sprite_type(1), B => L2_n_474, ZN => L2_n_494);
  L2_g12491 : AOI22D0BWP7T port map(A1 => L2_n_484, A2 => L2_n_270, B1 => L2_n_431, B2 => L2_n_263, ZN => L2_n_493);
  L2_g12492 : AN2D0BWP7T port map(A1 => L2_n_487, A2 => L2_n_439, Z => L2_n_492);
  L2_g12493 : AO211D0BWP7T port map(A1 => L2_n_430, A2 => L2_n_267, B => L2_n_461, C => L2_n_462, Z => L2_n_546);
  L2_g12494 : OAI22D0BWP7T port map(A1 => L2_n_468, A2 => L2_n_272, B1 => L2_n_390, B2 => L2_n_312, ZN => L2_n_491);
  L2_g12495 : AOI31D0BWP7T port map(A1 => L2_n_450, A2 => L2_n_419, A3 => L2_n_270, B => L2_n_480, ZN => L2_n_490);
  L2_g12496 : OAI22D0BWP7T port map(A1 => L2_n_470, A2 => L2_n_223, B1 => L2_n_378, B2 => L2_n_265, ZN => L2_n_489);
  L2_g12497 : AOI221D0BWP7T port map(A1 => L2_n_239, A2 => L2_n_311, B1 => L2_n_243, B2 => L2_n_254, C => L2_n_463, ZN => L2_n_487);
  L2_g12498 : OAI21D0BWP7T port map(A1 => L2_n_447, A2 => L2_n_433, B => L2_n_263, ZN => L2_n_486);
  L2_g12499 : IND2D1BWP7T port map(A1 => L2_n_272, B1 => L2_n_465, ZN => L2_n_485);
  L2_g12500 : AOI211D1BWP7T port map(A1 => L2_n_330, A2 => L2_n_308, B => L2_n_442, C => L2_n_374, ZN => L2_n_484);
  L2_g12501 : ND4D0BWP7T port map(A1 => L2_n_450, A2 => L2_n_405, A3 => L2_n_409, A4 => L2_n_270, ZN => L2_n_483);
  L2_g12502 : AO221D0BWP7T port map(A1 => L2_n_406, A2 => L2_vgacontrol_vcount(8), B1 => L2_n_435, B2 => L2_vgacontrol_hcount(8), C => reset, Z => L2_n_482);
  L2_g12503 : OA21D0BWP7T port map(A1 => L2_n_289, A2 => L2_n_317, B => L2_n_472, Z => L2_n_481);
  L2_g12504 : NR4D0BWP7T port map(A1 => L2_n_432, A2 => L2_vgacontrol_hcount(1), A3 => L2_vgacontrol_hcount(0), A4 => L2_vgacontrol_hcount(3), ZN => L2_n_488);
  L2_g12505 : AOI211D1BWP7T port map(A1 => L2_n_421, A2 => L2_in_go_sprite_type(2), B => L2_n_459, C => L2_n_272, ZN => L2_n_480);
  L2_g12506 : OAI22D0BWP7T port map(A1 => L2_n_449, A2 => L2_n_223, B1 => L2_n_445, B2 => L2_n_250, ZN => L2_n_479);
  L2_g12507 : OAI22D0BWP7T port map(A1 => L2_n_458, A2 => L2_n_280, B1 => L2_n_349, B2 => L2_n_299, ZN => L2_n_478);
  L2_g12508 : OAI22D0BWP7T port map(A1 => L2_n_457, A2 => L2_n_280, B1 => L2_n_387, B2 => L2_score_score_sprite_type(1), ZN => L2_n_477);
  L2_g12509 : IND4D0BWP7T port map(A1 => L2_n_374, B1 => L2_n_295, B2 => L2_n_383, B3 => L2_n_418, ZN => L2_n_476);
  L2_g12510 : OA22D0BWP7T port map(A1 => L2_n_452, A2 => L2_n_277, B1 => L2_n_317, B2 => L2_n_365, Z => L2_n_475);
  L2_g12511 : MOAI22D0BWP7T port map(A1 => L2_n_309, A2 => L2_n_292, B1 => L2_n_451, B2 => L2_n_276, ZN => L2_n_474);
  L2_g12512 : MAOI22D0BWP7T port map(A1 => L2_n_441, A2 => L2_score_score_sprite_type(1), B1 => L2_n_293, B2 => L2_n_299, ZN => L2_n_473);
  L2_g12513 : OAI221D0BWP7T port map(A1 => L2_n_336, A2 => L2_n_257, B1 => L2_n_233, B2 => L2_n_286, C => L2_n_440, ZN => L2_n_470);
  L2_g12514 : AOI221D0BWP7T port map(A1 => L2_n_331, A2 => L2_n_315, B1 => L2_n_238, B2 => L2_n_313, C => L2_n_460, ZN => L2_n_469);
  L2_g12515 : NR2XD0BWP7T port map(A1 => L2_n_460, A2 => L2_n_366, ZN => L2_n_468);
  L2_g12516 : IIND4D0BWP7T port map(A1 => L2_n_438, A2 => L2_n_374, B1 => L2_n_392, B2 => L2_n_409, ZN => L2_n_467);
  L2_g12517 : OR2D1BWP7T port map(A1 => L2_n_453, A2 => L2_n_277, Z => L2_n_472);
  L2_g12518 : OAI21D0BWP7T port map(A1 => L2_n_414, A2 => L2_n_340, B => L2_n_276, ZN => L2_n_471);
  L2_g12519 : ND4D0BWP7T port map(A1 => L2_n_427, A2 => L2_n_381, A3 => L2_n_359, A4 => L2_n_270, ZN => L2_n_466);
  L2_g12520 : OAI31D0BWP7T port map(A1 => L2_in_go_sprite_type(0), A2 => L2_n_236, A3 => L2_n_369, B => L2_n_444, ZN => L2_n_465);
  L2_g12521 : AOI211XD0BWP7T port map(A1 => L2_n_362, A2 => L2_n_311, B => L2_n_422, C => L2_n_382, ZN => L2_n_464);
  L2_g12522 : OAI222D0BWP7T port map(A1 => L2_n_389, A2 => L2_score_score_sprite_type(2), B1 => L2_n_319, B2 => L2_n_329, C1 => L2_n_260, C2 => L2_n_346, ZN => L2_n_463);
  L2_g12523 : OAI22D0BWP7T port map(A1 => L2_n_434, A2 => L2_n_275, B1 => L2_n_345, B2 => L2_n_319, ZN => L2_n_462);
  L2_g12524 : OAI22D0BWP7T port map(A1 => L2_n_420, A2 => L2_n_280, B1 => L2_n_399, B2 => L2_n_277, ZN => L2_n_461);
  L2_g12525 : AOI211XD0BWP7T port map(A1 => L2_n_376, A2 => L2_in_go_sprite_type(1), B => L2_n_357, C => L2_n_250, ZN => L2_n_459);
  L2_g12526 : AOI211XD0BWP7T port map(A1 => L2_n_361, A2 => L2_n_258, B => L2_n_385, C => L2_n_412, ZN => L2_n_458);
  L2_g12527 : AOI211XD0BWP7T port map(A1 => L2_n_377, A2 => L2_n_235, B => L2_n_388, C => L2_n_412, ZN => L2_n_457);
  L2_g12528 : OAI221D0BWP7T port map(A1 => L2_n_296, A2 => L2_n_260, B1 => L2_n_259, B2 => L2_n_249, C => L2_n_426, ZN => L2_n_456);
  L2_g12529 : AOI31D0BWP7T port map(A1 => L2_n_303, A2 => L2_n_276, A3 => L2_n_259, B => L2_n_429, ZN => L2_n_455);
  L2_g12530 : AOI211XD0BWP7T port map(A1 => L2_n_344, A2 => L2_n_313, B => L2_n_417, C => L2_n_395, ZN => L2_n_454);
  L2_g12531 : AOI21D0BWP7T port map(A1 => L2_n_361, A2 => L2_n_235, B => L2_n_425, ZN => L2_n_453);
  L2_g12532 : AOI21D0BWP7T port map(A1 => L2_n_344, A2 => L2_n_235, B => L2_n_425, ZN => L2_n_452);
  L2_g12533 : OAI211D1BWP7T port map(A1 => L2_n_259, A2 => L2_n_307, B => L2_n_426, C => L2_n_368, ZN => L2_n_451);
  L2_g12534 : OAI211D1BWP7T port map(A1 => L2_n_252, A2 => L2_n_375, B => L2_n_396, C => L2_n_326, ZN => L2_n_460);
  L2_g12535 : OAI222D0BWP7T port map(A1 => L2_n_369, A2 => L2_n_257, B1 => L2_n_244, B2 => L2_n_365, C1 => L2_n_261, C2 => L2_n_309, ZN => L2_n_449);
  L2_g12536 : OAI22D0BWP7T port map(A1 => L2_n_400, A2 => L2_score_score_sprite_type(3), B1 => L2_n_278, B2 => L2_n_317, ZN => L2_n_448);
  L2_g12537 : OAI22D0BWP7T port map(A1 => L2_n_408, A2 => L2_n_269, B1 => L2_n_278, B2 => L2_n_295, ZN => L2_n_447);
  L2_g12538 : OAI211D1BWP7T port map(A1 => L2_n_386, A2 => L2_n_380, B => L2_n_263, C => L2_n_223, ZN => L2_n_446);
  L2_g12539 : OAI222D0BWP7T port map(A1 => L2_n_393, A2 => L2_n_227, B1 => L2_n_257, B2 => L2_n_325, C1 => L2_n_233, C2 => L2_n_279, ZN => L2_n_445);
  L2_g12540 : IAO21D0BWP7T port map(A1 => L2_n_393, A2 => L2_n_252, B => L2_n_401, ZN => L2_n_444);
  L2_g12541 : OA222D0BWP7T port map(A1 => L2_n_375, A2 => L2_n_227, B1 => L2_n_257, B2 => L2_n_345, C1 => L2_n_233, C2 => L2_n_320, Z => L2_n_443);
  L2_g12542 : OAI22D0BWP7T port map(A1 => L2_n_404, A2 => L2_n_353, B1 => L2_n_338, B2 => L2_n_269, ZN => L2_n_442);
  L2_g12543 : MOAI22D0BWP7T port map(A1 => L2_n_402, A2 => L2_score_score_sprite_type(2), B1 => L2_n_361, B2 => L2_n_311, ZN => L2_n_441);
  L2_g12544 : MAOI22D0BWP7T port map(A1 => L2_n_407, A2 => L2_in_go_sprite_type(1), B1 => L2_n_289, B2 => L2_n_261, ZN => L2_n_440);
  L2_g12545 : AOI31D0BWP7T port map(A1 => L2_n_362, A2 => L2_n_268, A3 => L2_in_go_sprite_type(0), B => L2_n_437, ZN => L2_n_450);
  L2_g12546 : OAI22D0BWP7T port map(A1 => L2_n_361, A2 => L2_n_337, B1 => L2_n_257, B2 => L2_n_223, ZN => L2_n_437);
  L2_g12547 : AOI31D0BWP7T port map(A1 => L2_n_321, A2 => L2_vgacontrol_vcount(7), A3 => L2_vgacontrol_vcount(8), B => L2_n_411, ZN => L2_n_436);
  L2_g12548 : OR3D1BWP7T port map(A1 => L2_vgacontrol_hcount(7), A2 => L2_vgacontrol_hcount(6), A3 => L2_n_371, Z => L2_n_435);
  L2_g12549 : AOI211XD0BWP7T port map(A1 => L2_n_353, A2 => L2_score_score_sprite_type(3), B => L2_n_347, C => L2_n_290, ZN => L2_n_434);
  L2_g12550 : MOAI22D0BWP7T port map(A1 => L2_n_372, A2 => L2_n_236, B1 => L2_n_378, B2 => L2_n_264, ZN => L2_n_433);
  L2_g12551 : IIND4D0BWP7T port map(A1 => L2_vgacontrol_hcount(7), A2 => L2_vgacontrol_hcount(8), B1 => L2_n_322, B2 => L2_vgacontrol_hcount(6), ZN => L2_n_432);
  L2_g12552 : OAI22D0BWP7T port map(A1 => L2_n_370, A2 => L2_n_265, B1 => L2_n_364, B2 => L2_n_252, ZN => L2_n_431);
  L2_g12553 : AO21D0BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_n_258, B => L2_n_394, Z => L2_n_430);
  L2_g12554 : AOI211D0BWP7T port map(A1 => L2_n_348, A2 => L2_n_278, B => L2_n_266, C => L2_score_score_sprite_type(3), ZN => L2_n_429);
  L2_g12555 : AOI31D0BWP7T port map(A1 => L2_n_318, A2 => L2_in_go_sprite_type(0), A3 => L2_in_go_sprite_type(2), B => L2_n_391, ZN => L2_n_428);
  L2_g12556 : OAI21D0BWP7T port map(A1 => L2_n_362, A2 => L2_in_go_sprite_type(2), B => L2_n_256, ZN => L2_n_427);
  L2_g12557 : IOA21D1BWP7T port map(A1 => L2_n_373, A2 => L2_n_260, B => L2_score_score_sprite_type(2), ZN => L2_n_439);
  L2_g12558 : NR2XD0BWP7T port map(A1 => L2_n_407, A2 => L2_n_269, ZN => L2_n_438);
  L2_g12559 : OA222D0BWP7T port map(A1 => L2_n_376, A2 => L2_n_227, B1 => L2_n_257, B2 => L2_n_340, C1 => L2_n_233, C2 => L2_n_287, Z => L2_n_423);
  L2_g12560 : AO32D1BWP7T port map(A1 => L2_n_291, A2 => L2_n_235, A3 => L2_n_225, B1 => L2_n_360, B2 => L2_n_254, Z => L2_n_422);
  L2_g12561 : OA222D0BWP7T port map(A1 => L2_n_349, A2 => L2_n_244, B1 => L2_n_261, B2 => L2_n_304, C1 => L2_n_257, C2 => L2_n_273, Z => L2_n_421);
  L2_g12562 : OA21D0BWP7T port map(A1 => L2_n_364, A2 => L2_score_score_sprite_type(3), B => L2_n_398, Z => L2_n_420);
  L2_g12563 : AOI222D0BWP7T port map(A1 => L2_n_352, A2 => L2_n_284, B1 => L2_n_341, B2 => L2_n_308, C1 => L2_n_293, C2 => L2_n_237, ZN => L2_n_419);
  L2_g12564 : AOI22D0BWP7T port map(A1 => L2_n_362, A2 => L2_n_315, B1 => L2_n_327, B2 => L2_n_223, ZN => L2_n_418);
  L2_g12565 : OAI22D0BWP7T port map(A1 => L2_n_365, A2 => L2_n_295, B1 => L2_n_278, B2 => L2_n_236, ZN => L2_n_417);
  L2_g12566 : OA21D0BWP7T port map(A1 => L2_n_300, A2 => L2_n_233, B => L2_n_379, Z => L2_n_416);
  L2_g12567 : AOI22D0BWP7T port map(A1 => L2_n_377, A2 => L2_n_335, B1 => L2_n_242, B2 => L2_n_351, ZN => L2_n_415);
  L2_g12568 : AOI22D0BWP7T port map(A1 => L2_n_360, A2 => L2_score_score_sprite_type(3), B1 => L2_n_350, B2 => L2_n_228, ZN => L2_n_414);
  L2_g12569 : MAOI22D0BWP7T port map(A1 => L2_n_361, A2 => L2_n_351, B1 => L2_n_352, B2 => L2_n_334, ZN => L2_n_413);
  L2_g12570 : AOI22D0BWP7T port map(A1 => L2_n_363, A2 => L2_n_248, B1 => L2_n_329, B2 => L2_n_235, ZN => L2_n_426);
  L2_g12571 : OAI22D0BWP7T port map(A1 => L2_n_360, A2 => L2_n_247, B1 => L2_n_243, B2 => L2_n_260, ZN => L2_n_425);
  L2_g12572 : IND4D0BWP7T port map(A1 => L2_n_250, B1 => L2_in_go_sprite_type(3), B2 => L2_n_256, B3 => L2_n_355, ZN => L2_n_424);
  L2_g12573 : INVD0BWP7T port map(I => L2_n_407, ZN => L2_n_408);
  L2_g12574 : NR2D1BWP7T port map(A1 => L2_n_358, A2 => L2_n_522, ZN => L2_n_406);
  L2_g12575 : AOI22D0BWP7T port map(A1 => L2_n_333, A2 => L2_n_284, B1 => L2_n_349, B2 => L2_n_237, ZN => L2_n_405);
  L2_g12576 : IAO21D0BWP7T port map(A1 => L2_n_338, A2 => L2_n_265, B => L2_n_284, ZN => L2_n_404);
  L2_g12577 : AO21D0BWP7T port map(A1 => L2_n_306, A2 => L2_n_316, B => L2_n_366, Z => L2_n_403);
  L2_g12578 : OA21D0BWP7T port map(A1 => L2_n_352, A2 => L2_score_score_sprite_type(0), B => L2_n_341, Z => L2_n_402);
  L2_g12579 : AOI21D0BWP7T port map(A1 => L2_n_339, A2 => L2_n_279, B => L2_n_265, ZN => L2_n_401);
  L2_g12580 : AO21D0BWP7T port map(A1 => L2_n_348, A2 => L2_n_286, B => L2_n_266, Z => L2_n_400);
  L2_g12581 : AOI211XD0BWP7T port map(A1 => L2_n_242, A2 => L2_score_score_sprite_type(3), B => L2_n_342, C => L2_n_347, ZN => L2_n_399);
  L2_g12582 : AOI21D0BWP7T port map(A1 => L2_n_353, A2 => L2_n_248, B => L2_n_367, ZN => L2_n_398);
  L2_g12583 : OAI21D0BWP7T port map(A1 => L2_n_338, A2 => L2_n_314, B => L2_n_298, ZN => L2_n_397);
  L2_g12584 : OAI211D1BWP7T port map(A1 => L2_n_241, A2 => L2_n_301, B => L2_n_237, C => L2_n_224, ZN => L2_n_396);
  L2_g12585 : AOI21D0BWP7T port map(A1 => L2_n_339, A2 => L2_n_307, B => L2_in_go_sprite_type(1), ZN => L2_n_395);
  L2_g12586 : NR2D1BWP7T port map(A1 => L2_n_364, A2 => L2_n_260, ZN => L2_n_412);
  L2_g12587 : NR4D0BWP7T port map(A1 => L2_n_321, A2 => L2_vgacontrol_vcount(9), A3 => L2_vgacontrol_vcount(7), A4 => L2_vgacontrol_vcount(8), ZN => L2_n_411);
  L2_g12588 : NR3D0BWP7T port map(A1 => L2_n_343, A2 => L2_n_312, A3 => L2_n_261, ZN => L2_n_410);
  L2_g12589 : ND2D1BWP7T port map(A1 => L2_n_364, A2 => L2_n_308, ZN => L2_n_409);
  L2_g12590 : NR2XD0BWP7T port map(A1 => L2_n_360, A2 => L2_in_go_sprite_type(0), ZN => L2_n_407);
  L2_g12591 : OA22D0BWP7T port map(A1 => L2_n_344, A2 => L2_n_285, B1 => L2_n_265, B2 => L2_n_303, Z => L2_n_392);
  L2_g12592 : AO22D0BWP7T port map(A1 => L2_n_349, A2 => L2_n_313, B1 => L2_n_237, B2 => L2_n_273, Z => L2_n_391);
  L2_g12593 : OA221D0BWP7T port map(A1 => L2_n_330, A2 => L2_n_244, B1 => L2_n_257, B2 => L2_n_246, C => L2_n_328, Z => L2_n_390);
  L2_g12594 : AOI22D0BWP7T port map(A1 => L2_n_354, A2 => L2_n_235, B1 => L2_n_296, B2 => L2_n_248, ZN => L2_n_389);
  L2_g12595 : MOAI22D0BWP7T port map(A1 => L2_n_243, A2 => L2_n_259, B1 => L2_n_344, B2 => L2_n_248, ZN => L2_n_388);
  L2_g12596 : MOAI22D0BWP7T port map(A1 => L2_n_282, A2 => L2_n_532, B1 => L2_screencontrol_n_58, B2 => L2_n_533, ZN => L2_user_reset_new);
  L2_g12597 : MAOI22D0BWP7T port map(A1 => L2_n_306, A2 => L2_n_311, B1 => L2_n_350, B2 => L2_n_255, ZN => L2_n_387);
  L2_g12598 : OAI22D0BWP7T port map(A1 => L2_n_354, A2 => L2_n_244, B1 => L2_n_239, B2 => L2_n_261, ZN => L2_n_386);
  L2_g12599 : OAI22D0BWP7T port map(A1 => L2_n_333, A2 => L2_n_247, B1 => L2_n_289, B2 => L2_n_234, ZN => L2_n_385);
  L2_g12600 : OA22D0BWP7T port map(A1 => L2_n_336, A2 => L2_n_292, B1 => L2_n_294, B2 => L2_n_286, Z => L2_n_384);
  L2_g12601 : MAOI22D0BWP7T port map(A1 => L2_n_243, A2 => L2_n_268, B1 => L2_n_346, B2 => L2_n_261, ZN => L2_n_383);
  L2_g12602 : OAI22D0BWP7T port map(A1 => L2_n_331, A2 => L2_n_323, B1 => L2_n_240, B2 => L2_n_260, ZN => L2_n_382);
  L2_g12603 : MAOI22D0BWP7T port map(A1 => L2_n_330, A2 => L2_n_316, B1 => L2_n_331, B2 => L2_n_285, ZN => L2_n_381);
  L2_g12604 : OAI22D0BWP7T port map(A1 => L2_n_330, A2 => L2_n_257, B1 => L2_n_249, B2 => L2_n_233, ZN => L2_n_380);
  L2_g12605 : MAOI22D0BWP7T port map(A1 => L2_n_331, A2 => L2_n_245, B1 => L2_n_309, B2 => L2_n_257, ZN => L2_n_379);
  L2_g12606 : MOAI22D0BWP7T port map(A1 => L2_n_350, A2 => L2_n_228, B1 => L2_n_241, B2 => L2_n_258, ZN => L2_n_394);
  L2_g12607 : AOI22D0BWP7T port map(A1 => L2_n_342, A2 => L2_in_go_sprite_type(0), B1 => L2_n_238, B2 => L2_n_224, ZN => L2_n_393);
  L2_g12609 : ND2D1BWP7T port map(A1 => L2_n_343, A2 => L2_score_score_sprite_type(0), ZN => L2_n_373);
  L2_g12610 : INR2XD0BWP7T port map(A1 => L2_n_286, B1 => L2_n_338, ZN => L2_n_372);
  L2_g12611 : NR2D0BWP7T port map(A1 => L2_n_526, A2 => L2_n_524, ZN => L2_n_371);
  L2_g12612 : NR2XD0BWP7T port map(A1 => L2_n_338, A2 => L2_n_290, ZN => L2_n_370);
  L2_g12613 : CKND2D1BWP7T port map(A1 => L2_n_332, A2 => L2_n_341, ZN => L2_n_378);
  L2_g12614 : IND2D1BWP7T port map(A1 => L2_n_238, B1 => L2_n_333, ZN => L2_n_377);
  L2_g12615 : IND2D1BWP7T port map(A1 => L2_n_355, B1 => L2_n_332, ZN => L2_n_376);
  L2_g12616 : NR2XD0BWP7T port map(A1 => L2_n_342, A2 => L2_n_338, ZN => L2_n_375);
  L2_g12617 : AN2D1BWP7T port map(A1 => L2_n_332, A2 => L2_n_237, Z => L2_n_374);
  L2_g12618 : INVD0BWP7T port map(I => L2_n_367, ZN => L2_n_368);
  L2_g12619 : INVD0BWP7T port map(I => L2_n_363, ZN => L2_n_362);
  L2_g12620 : INVD1BWP7T port map(I => L2_n_361, ZN => L2_n_360);
  L2_g12621 : AOI22D0BWP7T port map(A1 => L2_n_239, A2 => L2_n_308, B1 => L2_n_229, B2 => L2_n_237, ZN => L2_n_359);
  L2_g12622 : AOI21D0BWP7T port map(A1 => L2_n_302, A2 => L2_vgacontrol_vcount(4), B => L2_vgacontrol_vcount(5), ZN => L2_n_358);
  L2_g12623 : AO21D0BWP7T port map(A1 => L2_n_287, A2 => L2_n_232, B => L2_n_324, Z => L2_n_357);
  L2_g12624 : NR2XD0BWP7T port map(A1 => L2_n_329, A2 => L2_n_241, ZN => L2_n_369);
  L2_g12625 : NR2D0BWP7T port map(A1 => L2_n_330, A2 => L2_n_260, ZN => L2_n_367);
  L2_g12626 : INR2D0BWP7T port map(A1 => L2_n_315, B1 => L2_n_330, ZN => L2_n_366);
  L2_g12627 : NR3D0BWP7T port map(A1 => L2_n_305, A2 => L2_n_238, A3 => L2_n_241, ZN => L2_n_365);
  L2_g12628 : NR3D0BWP7T port map(A1 => L2_n_310, A2 => L2_n_240, A3 => L2_n_274, ZN => L2_n_364);
  L2_g12629 : AOI21D0BWP7T port map(A1 => L2_n_288, A2 => L2_county(2), B => L2_n_279, ZN => L2_n_363);
  L2_g12630 : ND2D1BWP7T port map(A1 => L2_n_341, A2 => L2_n_304, ZN => L2_n_361);
  L2_g12631 : INVD0BWP7T port map(I => L2_n_533, ZN => L2_n_356);
  L2_g12632 : INVD0BWP7T port map(I => L2_n_347, ZN => L2_n_348);
  L2_g12633 : INVD0BWP7T port map(I => L2_n_346, ZN => L2_n_345);
  L2_g12634 : INVD1BWP7T port map(I => L2_n_343, ZN => L2_n_342);
  L2_g12635 : INVD0BWP7T port map(I => L2_n_341, ZN => L2_n_340);
  L2_g12636 : INVD1BWP7T port map(I => L2_n_339, ZN => L2_n_338);
  L2_g12637 : NR2XD0BWP7T port map(A1 => L2_n_313, A2 => L2_n_264, ZN => L2_n_337);
  L2_g12638 : ND2D1BWP7T port map(A1 => L2_n_318, A2 => L2_n_304, ZN => L2_n_355);
  L2_g12639 : NR2D1BWP7T port map(A1 => L2_n_314, A2 => L2_n_306, ZN => L2_n_354);
  L2_g12640 : ND2D1BWP7T port map(A1 => L2_n_320, A2 => L2_n_253, ZN => L2_n_353);
  L2_g12641 : CKAN2D1BWP7T port map(A1 => L2_n_293, A2 => L2_n_281, Z => L2_n_352);
  L2_g12642 : AN2D1BWP7T port map(A1 => L2_n_308, A2 => L2_n_263, Z => L2_n_351);
  L2_g12643 : ND2D1BWP7T port map(A1 => L2_n_303, A2 => L2_score_score_sprite_type(0), ZN => L2_n_350);
  L2_g12644 : NR2XD0BWP7T port map(A1 => L2_n_305, A2 => L2_n_310, ZN => L2_n_349);
  L2_g12645 : INR2D1BWP7T port map(A1 => L2_n_303, B1 => L2_score_score_sprite_type(0), ZN => L2_n_347);
  L2_g12646 : ND2D1BWP7T port map(A1 => L2_n_318, A2 => L2_n_246, ZN => L2_n_346);
  L2_g12647 : ND2D1BWP7T port map(A1 => L2_n_288, A2 => L2_n_230, ZN => L2_n_344);
  L2_g12648 : NR2XD0BWP7T port map(A1 => L2_n_314, A2 => L2_n_310, ZN => L2_n_343);
  L2_g12649 : NR2XD0BWP7T port map(A1 => L2_n_310, A2 => L2_n_306, ZN => L2_n_341);
  L2_g12650 : ND2D1BWP7T port map(A1 => L2_n_303, A2 => L2_n_224, ZN => L2_n_339);
  L2_g12651 : INVD0BWP7T port map(I => L2_n_334, ZN => L2_n_335);
  L2_g12652 : INVD1BWP7T port map(I => L2_n_330, ZN => L2_n_329);
  L2_g12653 : OAI21D0BWP7T port map(A1 => L2_n_240, A2 => L2_n_241, B => L2_n_232, ZN => L2_n_328);
  L2_g12654 : OA21D0BWP7T port map(A1 => L2_n_232, A2 => L2_n_245, B => L2_n_296, Z => L2_n_327);
  L2_g12655 : IOA21D1BWP7T port map(A1 => L2_n_249, A2 => L2_n_230, B => L2_n_316, ZN => L2_n_326);
  L2_g12656 : NR2XD0BWP7T port map(A1 => L2_n_287, A2 => L2_n_274, ZN => L2_n_325);
  L2_g12657 : AOI21D0BWP7T port map(A1 => L2_n_251, A2 => L2_n_281, B => L2_n_257, ZN => L2_n_324);
  L2_g12658 : OA21D0BWP7T port map(A1 => L2_n_247, A2 => L2_score_score_sprite_type(2), B => L2_n_319, Z => L2_n_323);
  L2_g12659 : NR4D0BWP7T port map(A1 => L2_vgacontrol_hcount(9), A2 => L2_vgacontrol_hcount(2), A3 => L2_vgacontrol_hcount(4), A4 => L2_vgacontrol_hcount(5), ZN => L2_n_322);
  L2_g12660 : ND3D0BWP7T port map(A1 => L2_n_527, A2 => L2_vgacontrol_hcount(3), A3 => L2_vgacontrol_hcount(2), ZN => L2_n_526);
  L2_g12661 : INR2D1BWP7T port map(A1 => L2_n_309, B1 => L2_n_238, ZN => L2_n_336);
  L2_g12662 : ND2D1BWP7T port map(A1 => L2_n_284, A2 => L2_n_263, ZN => L2_n_334);
  L2_g12663 : CKAN2D1BWP7T port map(A1 => L2_n_286, A2 => L2_n_304, Z => L2_n_333);
  L2_g12664 : ND2D1BWP7T port map(A1 => L2_n_303, A2 => L2_in_go_sprite_type(0), ZN => L2_n_332);
  L2_g12665 : ND2D1BWP7T port map(A1 => L2_n_309, A2 => L2_n_239, ZN => L2_n_331);
  L2_g12666 : INR2XD0BWP7T port map(A1 => L2_n_253, B1 => L2_n_301, ZN => L2_n_330);
  L2_g12667 : INVD1BWP7T port map(I => L2_n_307, ZN => L2_n_306);
  L2_g12668 : INVD1BWP7T port map(I => L2_n_305, ZN => L2_n_304);
  L2_g12669 : OR2D1BWP7T port map(A1 => L2_n_529, A2 => L2_vgacontrol_vcount(6), Z => L2_n_321);
  L2_g12670 : NR2XD0BWP7T port map(A1 => L2_n_241, A2 => L2_in_go_y_pos(1), ZN => L2_n_320);
  L2_g12671 : ND2D1BWP7T port map(A1 => L2_n_235, A2 => L2_score_score_sprite_type(2), ZN => L2_n_319);
  L2_g12672 : IND2D1BWP7T port map(A1 => L2_n_249, B1 => L2_n_230, ZN => L2_n_318);
  L2_g12673 : OR2D1BWP7T port map(A1 => L2_n_277, A2 => L2_n_259, Z => L2_n_317);
  L2_g12674 : NR2D0BWP7T port map(A1 => L2_n_233, A2 => L2_in_go_sprite_type(2), ZN => L2_n_316);
  L2_g12675 : NR2D1BWP7T port map(A1 => L2_n_257, A2 => L2_in_go_sprite_type(2), ZN => L2_n_315);
  L2_g12676 : INR2D1BWP7T port map(A1 => L2_n_238, B1 => L2_county(0), ZN => L2_n_314);
  L2_g12677 : NR2D1BWP7T port map(A1 => L2_n_269, A2 => L2_in_go_sprite_type(0), ZN => L2_n_313);
  L2_g12678 : CKND2D1BWP7T port map(A1 => L2_n_263, A2 => L2_in_go_sprite_type(2), ZN => L2_n_312);
  L2_g12679 : NR2XD0BWP7T port map(A1 => L2_n_259, A2 => L2_score_score_sprite_type(2), ZN => L2_n_311);
  L2_g12680 : AN2D1BWP7T port map(A1 => L2_n_241, A2 => L2_n_229, Z => L2_n_310);
  L2_g12681 : IND2D1BWP7T port map(A1 => L2_n_246, B1 => L2_county(0), ZN => L2_n_309);
  L2_g12682 : NR2XD0BWP7T port map(A1 => L2_n_261, A2 => L2_in_go_sprite_type(2), ZN => L2_n_308);
  L2_g12683 : ND2D1BWP7T port map(A1 => L2_n_274, A2 => L2_county(0), ZN => L2_n_307);
  L2_g12684 : NR2XD0BWP7T port map(A1 => L2_n_246, A2 => L2_county(0), ZN => L2_n_305);
  L2_g12685 : ND2D1BWP7T port map(A1 => L2_n_243, A2 => L2_n_230, ZN => L2_n_303);
  L2_g12686 : INVD0BWP7T port map(I => L2_n_521, ZN => L2_n_302);
  L2_g12687 : CKND1BWP7T port map(I => L2_n_298, ZN => L2_n_297);
  L2_g12688 : INVD0BWP7T port map(I => L2_n_290, ZN => L2_n_291);
  L2_g12689 : INVD0BWP7T port map(I => L2_n_288, ZN => L2_n_287);
  L2_g12690 : INVD1BWP7T port map(I => L2_n_285, ZN => L2_n_284);
  L2_g12691 : NR3D0BWP7T port map(A1 => L2_n_530, A2 => L2_shift_L12_count_internal(1), A3 => L2_shift_L12_count_internal(0), ZN => L2_n_283);
  L2_g12692 : IND3D1BWP7T port map(A1 => L2_n_525, B1 => L2_vgacontrol_vcount(2), B2 => L2_vgacontrol_vcount(3), ZN => L2_n_521);
  L2_g12693 : IND2D1BWP7T port map(A1 => L2_n_238, B1 => L2_n_246, ZN => L2_n_301);
  L2_g12694 : AN2D0BWP7T port map(A1 => L2_n_253, A2 => L2_n_251, Z => L2_n_300);
  L2_g12695 : IND2D1BWP7T port map(A1 => L2_n_260, B1 => L2_n_267, ZN => L2_n_299);
  L2_g12696 : NR2D0BWP7T port map(A1 => L2_n_272, A2 => L2_n_269, ZN => L2_n_298);
  L2_g12697 : NR2D1BWP7T port map(A1 => L2_n_238, A2 => L2_n_240, ZN => L2_n_296);
  L2_g12698 : OR2D1BWP7T port map(A1 => L2_n_261, A2 => L2_n_223, Z => L2_n_295);
  L2_g12699 : ND2D1BWP7T port map(A1 => L2_n_267, A2 => L2_n_258, ZN => L2_n_294);
  L2_g12700 : CKAN2D1BWP7T port map(A1 => L2_n_251, A2 => L2_n_246, Z => L2_n_293);
  L2_g12701 : ND2D1BWP7T port map(A1 => L2_n_267, A2 => L2_n_235, ZN => L2_n_292);
  L2_g12702 : IND2D1BWP7T port map(A1 => L2_n_238, B1 => L2_n_249, ZN => L2_n_290);
  L2_g12703 : AN2D1BWP7T port map(A1 => L2_n_251, A2 => L2_n_273, Z => L2_n_289);
  L2_g12704 : CKND2D1BWP7T port map(A1 => L2_n_249, A2 => L2_n_242, ZN => L2_n_288);
  L2_g12705 : INR2D1BWP7T port map(A1 => L2_n_249, B1 => L2_n_241, ZN => L2_n_286);
  L2_g12706 : ND2D1BWP7T port map(A1 => L2_n_245, A2 => L2_n_223, ZN => L2_n_285);
  L2_g12707 : MOAI22D0BWP7T port map(A1 => L2_screencontrol_state(1), A2 => L2_screencontrol_state(0), B1 => L2_screencontrol_state(0), B2 => L2_screencontrol_state(1), ZN => L2_n_533);
  L2_g12708 : INVD0BWP7T port map(I => L2_n_282, ZN => L2_screencontrol_n_66);
  L2_g12709 : INVD0BWP7T port map(I => L2_n_276, ZN => L2_n_275);
  L2_g12710 : INVD0BWP7T port map(I => L2_n_274, ZN => L2_n_273);
  L2_g12711 : INVD1BWP7T port map(I => L2_n_271, ZN => L2_n_270);
  L2_g12712 : INVD0BWP7T port map(I => L2_n_269, ZN => L2_n_268);
  L2_g12713 : INVD0BWP7T port map(I => L2_n_267, ZN => L2_n_266);
  L2_g12714 : INVD0BWP7T port map(I => L2_n_265, ZN => L2_n_264);
  L2_g12715 : INVD0BWP7T port map(I => L2_n_263, ZN => L2_n_262);
  L2_g12716 : INVD1BWP7T port map(I => L2_n_259, ZN => L2_n_258);
  L2_g12717 : INVD0BWP7T port map(I => L2_n_257, ZN => L2_n_256);
  L2_g12718 : CKAN2D1BWP7T port map(A1 => L2_vgacontrol_vcount(4), A2 => L2_vgacontrol_vcount(5), Z => L2_n_529);
  L2_g12719 : ND2D1BWP7T port map(A1 => L2_calc_start_internal, A2 => L2_screencontrol_go, ZN => L2_n_282);
  L2_g12720 : IND2D1BWP7T port map(A1 => L2_shift_shift_clock_reset, B1 => L2_shift_L12_count_internal(2), ZN => L2_n_530);
  L2_g12721 : CKND2D1BWP7T port map(A1 => L2_vgacontrol_vcount(1), A2 => L2_vgacontrol_vcount(0), ZN => L2_n_525);
  L2_g12722 : CKND2D0BWP7T port map(A1 => L2_county(0), A2 => L2_county(2), ZN => L2_n_281);
  L2_g12723 : ND2D1BWP7T port map(A1 => L2_n_225, A2 => L2_score_score_sprite_type(1), ZN => L2_n_280);
  L2_g12724 : NR2XD0BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(2), ZN => L2_n_279);
  L2_g12725 : NR2XD0BWP7T port map(A1 => L2_county(2), A2 => L2_county(0), ZN => L2_n_278);
  L2_g12726 : ND2D1BWP7T port map(A1 => L2_score_score_sprite_type(2), A2 => L2_score_score_sprite_type(1), ZN => L2_n_277);
  L2_g12727 : NR2D0BWP7T port map(A1 => L2_score_score_sprite_type(2), A2 => L2_score_score_sprite_type(1), ZN => L2_n_276);
  L2_g12728 : NR2XD0BWP7T port map(A1 => L2_n_229, A2 => L2_n_230, ZN => L2_n_274);
  L2_g12729 : IND2D1BWP7T port map(A1 => L2_in_go_sprite_type(3), B1 => L2_in_go_sprite_type(4), ZN => L2_n_272);
  L2_g12730 : CKND2D1BWP7T port map(A1 => L2_n_231, A2 => L2_in_go_sprite_type(3), ZN => L2_n_271);
  L2_g12731 : ND2D1BWP7T port map(A1 => L2_in_go_sprite_type(1), A2 => L2_in_go_sprite_type(2), ZN => L2_n_269);
  L2_g12732 : NR2D1BWP7T port map(A1 => L2_n_225, A2 => L2_score_score_sprite_type(1), ZN => L2_n_267);
  L2_g12733 : ND2D1BWP7T port map(A1 => L2_n_223, A2 => L2_n_227, ZN => L2_n_265);
  L2_g12734 : NR2D1BWP7T port map(A1 => L2_in_go_sprite_type(3), A2 => L2_in_go_sprite_type(4), ZN => L2_n_263);
  L2_g12735 : ND2D1BWP7T port map(A1 => L2_in_go_sprite_type(0), A2 => L2_in_go_sprite_type(1), ZN => L2_n_261);
  L2_g12736 : ND2D1BWP7T port map(A1 => L2_score_score_sprite_type(3), A2 => L2_score_score_sprite_type(0), ZN => L2_n_260);
  L2_g12737 : CKND2D1BWP7T port map(A1 => L2_n_228, A2 => L2_score_score_sprite_type(0), ZN => L2_n_259);
  L2_g12738 : ND2D1BWP7T port map(A1 => L2_n_227, A2 => L2_n_224, ZN => L2_n_257);
  L2_g12739 : INVD0BWP7T port map(I => L2_n_254, ZN => L2_n_255);
  L2_g12740 : INVD0BWP7T port map(I => L2_n_248, ZN => L2_n_247);
  L2_g12741 : INVD1BWP7T port map(I => L2_n_245, ZN => L2_n_244);
  L2_g12742 : INVD0BWP7T port map(I => L2_n_243, ZN => L2_n_242);
  L2_g12743 : INVD1BWP7T port map(I => L2_n_240, ZN => L2_n_239);
  L2_g12744 : INVD0BWP7T port map(I => L2_n_237, ZN => L2_n_236);
  L2_g12745 : INVD0BWP7T port map(I => L2_n_235, ZN => L2_n_234);
  L2_g12746 : INVD0BWP7T port map(I => L2_n_233, ZN => L2_n_232);
  L2_g12747 : NR2XD0BWP7T port map(A1 => L2_vgacontrol_vcount(5), A2 => L2_vgacontrol_vcount(6), ZN => L2_n_528);
  L2_g12748 : IND2D1BWP7T port map(A1 => L2_screencontrol_state(0), B1 => L2_screencontrol_state(1), ZN => L2_n_532);
  L2_g12749 : AN2D1BWP7T port map(A1 => L2_vgacontrol_hcount(0), A2 => L2_vgacontrol_hcount(1), Z => L2_n_527);
  L2_g12750 : CKND2D1BWP7T port map(A1 => L2_vgacontrol_hcount(4), A2 => L2_vgacontrol_hcount(5), ZN => L2_n_524);
  L2_g12751 : NR2XD0BWP7T port map(A1 => L2_n_228, A2 => L2_n_225, ZN => L2_n_254);
  L2_g12752 : CKND2D1BWP7T port map(A1 => L2_vgacontrol_vcount(7), A2 => L2_vgacontrol_vcount(6), ZN => L2_n_522);
  L2_g12753 : CKND2D1BWP7T port map(A1 => L2_n_226, A2 => L2_county(2), ZN => L2_n_253);
  L2_g12754 : CKND2D1BWP7T port map(A1 => L2_n_223, A2 => L2_in_go_sprite_type(1), ZN => L2_n_252);
  L2_g12755 : ND2D1BWP7T port map(A1 => L2_n_229, A2 => L2_county(0), ZN => L2_n_251);
  L2_g12756 : ND2D1BWP7T port map(A1 => L2_n_223, A2 => L2_in_go_sprite_type(4), ZN => L2_n_250);
  L2_g12757 : CKND2D1BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(0), ZN => L2_n_249);
  L2_g12758 : NR2D1BWP7T port map(A1 => L2_n_228, A2 => L2_score_score_sprite_type(0), ZN => L2_n_248);
  L2_g12759 : CKND2D1BWP7T port map(A1 => L2_n_229, A2 => L2_county(2), ZN => L2_n_246);
  L2_g12760 : NR2XD0BWP7T port map(A1 => L2_n_227, A2 => L2_in_go_sprite_type(0), ZN => L2_n_245);
  L2_g12761 : NR2XD0BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(0), ZN => L2_n_243);
  L2_g12762 : NR2D1BWP7T port map(A1 => L2_n_226, A2 => L2_county(2), ZN => L2_n_241);
  L2_g12763 : NR2D1BWP7T port map(A1 => L2_n_229, A2 => L2_county(0), ZN => L2_n_240);
  L2_g12764 : NR2D1BWP7T port map(A1 => L2_n_229, A2 => L2_county(2), ZN => L2_n_238);
  L2_g12765 : NR2D1BWP7T port map(A1 => L2_in_go_sprite_type(1), A2 => L2_n_223, ZN => L2_n_237);
  L2_g12766 : NR2XD0BWP7T port map(A1 => L2_score_score_sprite_type(0), A2 => L2_score_score_sprite_type(3), ZN => L2_n_235);
  L2_g12767 : CKND2D1BWP7T port map(A1 => L2_n_227, A2 => L2_in_go_sprite_type(0), ZN => L2_n_233);
  L2_g12768 : INVD0BWP7T port map(I => L2_in_go_sprite_type(4), ZN => L2_n_231);
  L2_g12771 : INVD1BWP7T port map(I => L2_score_score_sprite_type(3), ZN => L2_n_228);
  L2_g12772 : INVD1BWP7T port map(I => L2_in_go_sprite_type(1), ZN => L2_n_227);
  L2_g12773 : INVD1BWP7T port map(I => L2_n_523, ZN => L2_calc_start_internal);
  L2_g12775 : INVD1BWP7T port map(I => L2_score_score_sprite_type(2), ZN => L2_n_225);
  L2_g12776 : INVD1BWP7T port map(I => L2_in_go_sprite_type(0), ZN => L2_n_224);
  L2_g12777 : INVD1BWP7T port map(I => L2_in_go_sprite_type(2), ZN => L2_n_223);
  L2_g4943 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gg(3), A2 => L2_n_539, B1 => L2_shift_pixel_arr_out_shift_gr(3), B2 => L2_n_538, C1 => L2_shift_pixel_arr_out_shift_pacman(3), C2 => L2_n_534, Z => L2_pixel_array_shifted(3));
  L2_g4944 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gr(5), A2 => L2_n_538, B1 => L2_shift_pixel_arr_out_shift_pacman(5), B2 => L2_n_534, C1 => L2_shift_pixel_arr_out_shift_gg(5), C2 => L2_n_539, Z => L2_pixel_array_shifted(5));
  L2_g4945 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gr(7), A2 => L2_n_538, B1 => L2_shift_pixel_arr_out_shift_pacman(7), B2 => L2_n_534, C1 => L2_shift_pixel_arr_out_shift_gg(7), C2 => L2_n_539, Z => L2_pixel_array_shifted(7));
  L2_g4946 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gg(2), A2 => L2_n_539, B1 => L2_shift_pixel_arr_out_shift_gr(2), B2 => L2_n_538, C1 => L2_shift_pixel_arr_out_shift_pacman(2), C2 => L2_n_534, Z => L2_pixel_array_shifted(2));
  L2_g4947 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gg(4), A2 => L2_n_539, B1 => L2_shift_pixel_arr_out_shift_gr(4), B2 => L2_n_538, C1 => L2_shift_pixel_arr_out_shift_pacman(4), C2 => L2_n_534, Z => L2_pixel_array_shifted(4));
  L2_g4948 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gg(1), A2 => L2_n_539, B1 => L2_shift_pixel_arr_out_shift_gr(1), B2 => L2_n_538, C1 => L2_shift_pixel_arr_out_shift_pacman(1), C2 => L2_n_534, Z => L2_pixel_array_shifted(1));
  L2_g4949 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gg(6), A2 => L2_n_539, B1 => L2_shift_pixel_arr_out_shift_gr(6), B2 => L2_n_538, C1 => L2_shift_pixel_arr_out_shift_pacman(6), C2 => L2_n_534, Z => L2_pixel_array_shifted(6));
  L2_g4950 : AO222D0BWP7T port map(A1 => L2_shift_pixel_arr_out_shift_gg(0), A2 => L2_n_539, B1 => L2_shift_pixel_arr_out_shift_gr(0), B2 => L2_n_538, C1 => L2_shift_pixel_arr_out_shift_pacman(0), C2 => L2_n_534, Z => L2_pixel_array_shifted(0));
  L2_g6387 : OR3D1BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_n_222, A3 => L2_n_219, Z => L2_pixel_array_to_shift(3));
  L2_g6388 : AO211D0BWP7T port map(A1 => L2_n_220, A2 => L2_n_172, B => L2_n_221, C => L2_n_222, Z => L2_pixel_array_to_shift(4));
  L2_g6389 : IND3D1BWP7T port map(A1 => L2_n_221, B1 => L2_n_214, B2 => L2_n_218, ZN => L2_pixel_array_to_shift(5));
  L2_g6390 : OAI211D1BWP7T port map(A1 => L2_n_180, A2 => L2_n_212, B => L2_n_218, C => L2_n_213, ZN => L2_pixel_array_to_shift(2));
  L2_g6391 : OAI222D0BWP7T port map(A1 => L2_n_212, A2 => L2_n_183, B1 => L2_n_177, B2 => L2_n_217, C1 => L2_n_201, C2 => L2_n_199, ZN => L2_n_222);
  L2_g6392 : OAI211D1BWP7T port map(A1 => L2_n_180, A2 => L2_n_199, B => L2_n_215, C => L2_n_213, ZN => L2_pixel_array_to_shift(1));
  L2_g6393 : OAI31D0BWP7T port map(A1 => L2_shift_cell_state_out_shift_pacman(3), A2 => L2_n_178, A3 => L2_n_212, B => L2_n_200, ZN => L2_n_221);
  L2_g6394 : OAI211D1BWP7T port map(A1 => L2_n_181, A2 => L2_n_199, B => L2_n_215, C => L2_n_213, ZN => L2_pixel_array_to_shift(6));
  L2_g6395 : OAI32D0BWP7T port map(A1 => L2_n_170, A2 => L2_shift_cell_state_out_shift_pacman(5), A3 => L2_n_212, B1 => L2_n_171, B2 => L2_n_210, ZN => L2_n_220);
  L2_g6396 : OAI33D1BWP7T port map(A1 => L2_n_171, A2 => L2_n_173, A3 => L2_n_212, B1 => L2_shift_cell_state_out_shift_pacman(3), B2 => L2_n_178, B3 => L2_n_210, ZN => L2_n_219);
  L2_g6397 : OA221D0BWP7T port map(A1 => L2_n_208, A2 => L2_n_201, B1 => L2_n_190, B2 => L2_n_191, C => L2_n_216, Z => L2_n_218);
  L2_g6398 : AOI211XD0BWP7T port map(A1 => L2_n_202, A2 => L2_shift_cell_state_out_shift_pacman(4), B => L2_n_209, C => L2_n_207, ZN => L2_n_217);
  L2_g6399 : MAOI22D0BWP7T port map(A1 => L2_n_203, A2 => L2_n_190, B1 => L2_n_197, B2 => L2_n_183, ZN => L2_n_216);
  L2_g6400 : OA22D0BWP7T port map(A1 => L2_n_205, A2 => L2_n_177, B1 => L2_n_171, B2 => L2_n_211, Z => L2_n_214);
  L2_g6401 : MAOI22D0BWP7T port map(A1 => L2_n_204, A2 => L2_n_172, B1 => L2_n_206, B2 => L2_n_183, ZN => L2_n_215);
  L2_g6402 : CKAN2D1BWP7T port map(A1 => L2_n_211, A2 => L2_n_200, Z => L2_n_213);
  L2_g6403 : CKAN2D1BWP7T port map(A1 => L2_n_206, A2 => L2_n_192, Z => L2_n_212);
  L2_g6404 : OAI21D0BWP7T port map(A1 => L2_n_184, A2 => L2_n_182, B => L2_n_201, ZN => L2_sprite_colour(0));
  L2_g6405 : AOI21D0BWP7T port map(A1 => L2_n_192, A2 => L2_n_195, B => L2_shift_cell_state_out_shift_pacman(4), ZN => L2_n_209);
  L2_g6406 : IND3D1BWP7T port map(A1 => L2_shift_cell_state_out_shift_pacman(5), B1 => L2_n_172, B2 => L2_n_196, ZN => L2_n_211);
  L2_g6407 : INR2XD0BWP7T port map(A1 => L2_n_192, B1 => L2_n_202, ZN => L2_n_210);
  L2_g6408 : INVD0BWP7T port map(I => L2_n_207, ZN => L2_n_208);
  L2_g6409 : AOI32D1BWP7T port map(A1 => L2_n_186, A2 => L2_n_190, A3 => L2_shift_cell_state_out_shift_pacman(4), B1 => L2_n_196, B2 => L2_n_168, ZN => L2_n_205);
  L2_g6410 : MOAI22D0BWP7T port map(A1 => L2_n_197, A2 => L2_n_190, B1 => L2_n_196, B2 => L2_n_190, ZN => L2_n_204);
  L2_g6411 : OAI22D0BWP7T port map(A1 => L2_n_195, A2 => L2_n_183, B1 => L2_n_188, B2 => L2_n_173, ZN => L2_n_203);
  L2_g6412 : MOAI22D0BWP7T port map(A1 => L2_n_197, A2 => L2_n_189, B1 => L2_n_198, B2 => L2_n_187, ZN => L2_n_207);
  L2_g6413 : OA21D0BWP7T port map(A1 => L2_n_189, A2 => L2_n_187, B => L2_n_199, Z => L2_n_206);
  L2_g6414 : NR2D1BWP7T port map(A1 => L2_n_198, A2 => L2_n_187, ZN => L2_n_202);
  L2_g6415 : ND2D1BWP7T port map(A1 => L2_n_193, A2 => L2_shift_cell_state_out_shift_pacman(2), ZN => L2_n_201);
  L2_g6416 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(7), ZN => L2_n_200);
  L2_g6417 : OAI21D0BWP7T port map(A1 => L2_n_184, A2 => L2_n_183, B => L2_n_194, ZN => L2_sprite_colour(2));
  L2_g6418 : OAI31D1BWP7T port map(A1 => L2_shift_cell_state_out_shift_pacman(1), A2 => L2_n_179, A3 => L2_n_184, B => L2_n_182, ZN => L2_pixel_array_to_shift(7));
  L2_g6419 : CKAN2D1BWP7T port map(A1 => L2_n_195, A2 => L2_n_197, Z => L2_n_199);
  L2_g6420 : INVD0BWP7T port map(I => L2_n_196, ZN => L2_n_195);
  L2_g6421 : NR2D1BWP7T port map(A1 => L2_n_190, A2 => L2_n_188, ZN => L2_n_198);
  L2_g6422 : ND2D1BWP7T port map(A1 => L2_n_186, A2 => L2_n_188, ZN => L2_n_197);
  L2_g6423 : NR2D1BWP7T port map(A1 => L2_n_186, A2 => L2_n_188, ZN => L2_n_196);
  L2_g6424 : INVD0BWP7T port map(I => L2_n_193, ZN => L2_n_194);
  L2_g6425 : IOA21D1BWP7T port map(A1 => L2_n_183, A2 => L2_n_173, B => L2_n_188, ZN => L2_n_191);
  L2_g6426 : NR3D0BWP7T port map(A1 => L2_n_185, A2 => L2_n_179, A3 => L2_shift_cell_state_out_shift_pacman(1), ZN => L2_n_193);
  L2_g6427 : ND2D1BWP7T port map(A1 => L2_n_189, A2 => L2_n_187, ZN => L2_n_192);
  L2_g6428 : INVD0BWP7T port map(I => L2_n_190, ZN => L2_n_189);
  L2_g6429 : INR2D1BWP7T port map(A1 => L2_n_182, B1 => L2_n_185, ZN => L2_sprite_colour(1));
  L2_g6430 : AOI222D0BWP7T port map(A1 => L2_n_534, A2 => L2_shift_y_pos_out_shift_pacman(0), B1 => L2_n_539, B2 => L2_shift_y_pos_out_shift_gg(0), C1 => L2_n_538, C2 => L2_shift_y_pos_out_shift_gr(0), ZN => L2_n_190);
  L2_g6431 : INVD1BWP7T port map(I => L2_n_187, ZN => L2_n_186);
  L2_g6432 : AOI222D0BWP7T port map(A1 => L2_n_534, A2 => L2_shift_y_pos_out_shift_pacman(1), B1 => L2_n_539, B2 => L2_shift_y_pos_out_shift_gg(1), C1 => L2_n_538, C2 => L2_shift_y_pos_out_shift_gr(1), ZN => L2_n_188);
  L2_g6433 : AOI222D0BWP7T port map(A1 => L2_n_534, A2 => L2_shift_y_pos_out_shift_pacman(2), B1 => L2_n_539, B2 => L2_shift_y_pos_out_shift_gg(2), C1 => L2_n_538, C2 => L2_shift_y_pos_out_shift_gr(2), ZN => L2_n_187);
  L2_g6434 : INVD0BWP7T port map(I => L2_n_185, ZN => L2_n_184);
  L2_g6435 : AOI21D0BWP7T port map(A1 => L2_n_534, A2 => L2_n_531, B => L2_n_539, ZN => L2_n_185);
  L2_g6436 : OA21D0BWP7T port map(A1 => L2_shift_cell_state_out_shift_pacman(2), A2 => L2_n_169, B => L2_n_534, Z => L2_n_183);
  L2_g6437 : ND3D0BWP7T port map(A1 => L2_n_534, A2 => L2_shift_cell_state_out_shift_pacman(2), A3 => L2_shift_cell_state_out_shift_pacman(1), ZN => L2_n_182);
  L2_g6438 : CKAN2D1BWP7T port map(A1 => L2_n_178, A2 => L2_n_177, Z => L2_n_181);
  L2_g6439 : NR3D0BWP7T port map(A1 => L2_n_172, A2 => L2_n_176, A3 => L2_n_174, ZN => L2_n_539);
  L2_g6440 : INVD0BWP7T port map(I => L2_n_534, ZN => L2_n_179);
  L2_g6441 : OA21D0BWP7T port map(A1 => L2_n_173, A2 => L2_n_168, B => L2_n_177, Z => L2_n_180);
  L2_g6442 : OAI21D0BWP7T port map(A1 => L2_n_175, A2 => L2_n_176, B => L2_n_173, ZN => L2_n_534);
  L2_g6443 : ND2D1BWP7T port map(A1 => L2_n_172, A2 => L2_n_168, ZN => L2_n_178);
  L2_g6444 : INR2D1BWP7T port map(A1 => L2_n_176, B1 => L2_n_172, ZN => L2_n_538);
  L2_g6445 : ND2D1BWP7T port map(A1 => L2_n_172, A2 => L2_shift_cell_state_out_shift_pacman(3), ZN => L2_n_177);
  L2_g6446 : INR3D0BWP7T port map(A1 => L2_shift_cell_state_out_shift_gr(1), B1 => L2_shift_cell_state_out_shift_gr(2), B2 => L2_shift_cell_state_out_shift_gr(0), ZN => L2_n_176);
  L2_g6447 : INVD1BWP7T port map(I => L2_n_174, ZN => L2_n_175);
  L2_g6448 : INVD1BWP7T port map(I => L2_n_173, ZN => L2_n_172);
  L2_g6449 : IND3D1BWP7T port map(A1 => L2_shift_cell_state_out_shift_gg(2), B1 => L2_shift_cell_state_out_shift_gg(1), B2 => L2_shift_cell_state_out_shift_gg(0), ZN => L2_n_174);
  L2_g6450 : IND3D1BWP7T port map(A1 => L2_shift_cell_state_out_shift_pacman(2), B1 => L2_n_169, B2 => L2_n_531, ZN => L2_n_173);
  L2_g6451 : ND2D1BWP7T port map(A1 => L2_n_170, A2 => L2_shift_cell_state_out_shift_pacman(4), ZN => L2_n_171);
  L2_g6452 : INVD0BWP7T port map(I => L2_shift_cell_state_out_shift_pacman(3), ZN => L2_n_170);
  L2_g6453 : INVD1BWP7T port map(I => L2_shift_cell_state_out_shift_pacman(1), ZN => L2_n_169);
  L2_g6454 : INVD1BWP7T port map(I => L2_shift_cell_state_out_shift_pacman(4), ZN => L2_n_168);
  L2_cnt_in_current_block_horizontal_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_46, D => L2_n_92, Q => L2_current_block_horizontal(0));
  L2_cnt_in_current_block_horizontal_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_46, D => L2_n_115, Q => L2_current_block_horizontal(1));
  L2_cnt_in_current_block_horizontal_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_46, D => L2_n_129, Q => L2_current_block_horizontal(2));
  L2_cnt_in_current_block_horizontal_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_46, D => L2_n_155, Q => L2_current_block_horizontal(3));
  L2_cnt_in_current_block_horizontal_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_46, D => L2_n_166, Q => L2_current_block_horizontal(4));
  L2_cnt_in_current_block_vertical_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_13, D => L2_n_35, Q => L2_current_block_vertical(0));
  L2_cnt_in_current_block_vertical_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_13, D => L2_n_101, Q => L2_current_block_vertical(1));
  L2_cnt_in_current_block_vertical_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_13, D => L2_n_119, Q => L2_current_block_vertical(2));
  L2_cnt_in_current_block_vertical_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_13, D => L2_n_136, Q => L2_current_block_vertical(3));
  L2_cnt_in_current_block_vertical_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_13, D => L2_n_163, Q => L2_current_block_vertical(4));
  L2_cnt_in_dual_pixel_y_reg : DFXQD1BWP7T port map(CP => clk, DA => L2_dual_pixel_y, DB => L2_n_41, SA => L2_n_71, Q => L2_dual_pixel_y);
  L2_screencontrol_go_reg : DFQD1BWP7T port map(CP => clk, D => L2_n_98, Q => L2_screencontrol_go);
  L2_screencontrol_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_n_110, Q => L2_screencontrol_state(0));
  L2_shift_L12_count_internal_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_n_116, Q => L2_shift_L12_count_internal(2));
  L2_shift_L13_current_pos_x_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_n_77, Q => L2_shift_pacman_pos_x(0));
  L2_shift_L13_current_pos_x_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_n_85, Q => L2_shift_pacman_pos_x(1));
  L2_shift_L13_current_pos_x_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_n_75, Q => L2_shift_pacman_pos_x(2));
  L2_shift_L13_current_pos_x_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_n_74, Q => L2_shift_pacman_pos_x(3));
  L2_shift_L13_current_pos_x_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_n_73, Q => L2_shift_pacman_pos_x(4));
  L2_shift_L13_current_pos_y_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_n_72, Q => L2_shift_pacman_pos_y(0));
  L2_shift_L13_current_pos_y_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_n_80, Q => L2_shift_pacman_pos_y(1));
  L2_shift_L13_current_pos_y_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_n_81, Q => L2_shift_pacman_pos_y(2));
  L2_shift_L13_current_pos_y_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_n_82, Q => L2_shift_pacman_pos_y(3));
  L2_shift_L13_current_pos_y_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_n_83, Q => L2_shift_pacman_pos_y(4));
  L2_shift_L22_current_pos_x_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_n_84, Q => L2_shift_gr_pos_x(0));
  L2_shift_L22_current_pos_x_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_n_70, Q => L2_shift_gr_pos_x(1));
  L2_shift_L22_current_pos_x_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_n_69, Q => L2_shift_gr_pos_x(2));
  L2_shift_L22_current_pos_x_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_n_68, Q => L2_shift_gr_pos_x(3));
  L2_shift_L22_current_pos_x_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_n_67, Q => L2_shift_gr_pos_x(4));
  L2_shift_L22_current_pos_y_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_n_66, Q => L2_shift_gr_pos_y(0));
  L2_shift_L22_current_pos_y_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_n_65, Q => L2_shift_gr_pos_y(1));
  L2_shift_L22_current_pos_y_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_n_64, Q => L2_shift_gr_pos_y(2));
  L2_shift_L22_current_pos_y_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_n_63, Q => L2_shift_gr_pos_y(3));
  L2_shift_L22_current_pos_y_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_n_62, Q => L2_shift_gr_pos_y(4));
  L2_shift_L32_current_pos_x_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_n_61, Q => L2_shift_gg_pos_x(0));
  L2_shift_L32_current_pos_x_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_n_60, Q => L2_shift_gg_pos_x(1));
  L2_shift_L32_current_pos_x_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_n_59, Q => L2_shift_gg_pos_x(2));
  L2_shift_L32_current_pos_x_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_n_58, Q => L2_shift_gg_pos_x(3));
  L2_shift_L32_current_pos_x_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_n_57, Q => L2_shift_gg_pos_x(4));
  L2_shift_L32_current_pos_y_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_n_56, Q => L2_shift_gg_pos_y(0));
  L2_shift_L32_current_pos_y_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_n_55, Q => L2_shift_gg_pos_y(1));
  L2_shift_L32_current_pos_y_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_n_54, Q => L2_shift_gg_pos_y(2));
  L2_shift_L32_current_pos_y_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_n_53, Q => L2_shift_gg_pos_y(3));
  L2_shift_L32_current_pos_y_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_n_52, Q => L2_shift_gg_pos_y(4));
  L2_vgacontrol_hcount_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_34, D => L2_n_117, Q => L2_vgacontrol_hcount(1));
  L2_vgacontrol_hcount_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_36, D => L2_n_117, Q => L2_vgacontrol_hcount(2));
  L2_vgacontrol_hcount_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_102, D => L2_n_117, Q => L2_vgacontrol_hcount(3));
  L2_vgacontrol_hcount_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_38, D => L2_n_117, Q => L2_vgacontrol_hcount(4));
  L2_vgacontrol_hcount_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_99, D => L2_n_117, Q => L2_vgacontrol_hcount(5));
  L2_vgacontrol_hcount_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_51, D => L2_n_117, Q => L2_vgacontrol_hcount(6));
  L2_vgacontrol_hcount_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_117, D => L2_n_107, Q => L2_vgacontrol_hcount(7));
  L2_vgacontrol_hcount_reg_8 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_117, D => L2_n_124, Q => L2_vgacontrol_hcount(8));
  L2_vgacontrol_hcount_reg_9 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_n_117, D => L2_n_145, Q => L2_vgacontrol_hcount(9));
  L2_vgacontrol_in_calc_start_game_reg : DFQD1BWP7T port map(CP => clk, D => L2_n_147, Q => calc_start_game_int);
  L2_vgacontrol_in_v_sync_reg : EDFKCNQD1BWP7T port map(CP => clk, CN => L2_n_2, D => L2_vgacontrol_vcount(1), E => L2_n_113, Q => L2_n_167);
  L2_vgacontrol_vcount_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_n_160, Q => L2_vgacontrol_vcount(1));
  L2_vgacontrol_vcount_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_n_162, Q => L2_vgacontrol_vcount(3));
  L2_vgacontrol_vcount_reg_5 : DFQD1BWP7T port map(CP => clk, D => L2_n_165, Q => L2_vgacontrol_vcount(5));
  L2_vgacontrol_vcount_reg_7 : DFQD1BWP7T port map(CP => clk, D => L2_n_164, Q => L2_vgacontrol_vcount(7));
  L2_vgacontrol_vcount_reg_8 : DFQD1BWP7T port map(CP => clk, D => L2_n_159, Q => L2_vgacontrol_vcount(8));
  L2_g7542 : MOAI22D0BWP7T port map(A1 => L2_n_154, A2 => L2_current_block_horizontal(4), B1 => L2_n_154, B2 => L2_current_block_horizontal(4), ZN => L2_n_166);
  L2_g7553 : AO21D0BWP7T port map(A1 => L2_n_149, A2 => L2_vgacontrol_vcount(5), B => L2_n_142, Z => L2_n_165);
  L2_g7554 : IOA21D1BWP7T port map(A1 => L2_n_148, A2 => L2_vgacontrol_vcount(7), B => L2_n_139, ZN => L2_n_164);
  L2_g7555 : MOAI22D0BWP7T port map(A1 => L2_n_135, A2 => L2_current_block_vertical(4), B1 => L2_n_135, B2 => L2_current_block_vertical(4), ZN => L2_n_163);
  L2_g7556 : IOA21D1BWP7T port map(A1 => L2_n_150, A2 => L2_vgacontrol_vcount(3), B => L2_n_161, ZN => L2_n_162);
  L2_g7559 : IND3D1BWP7T port map(A1 => L2_vgacontrol_vcount(3), B1 => L2_vgacontrol_vcount(2), B2 => L2_n_143, ZN => L2_n_161);
  L2_g7564 : OAI31D0BWP7T port map(A1 => L2_vgacontrol_vcount(1), A2 => L2_n_4, A3 => L2_n_134, B => L2_n_151, ZN => L2_n_160);
  L2_g7565 : OAI31D0BWP7T port map(A1 => L2_vgacontrol_vcount(8), A2 => L2_n_48, A3 => L2_n_134, B => L2_n_152, ZN => L2_n_159);
  L2_g7566 : OAI31D0BWP7T port map(A1 => L2_vgacontrol_vcount(6), A2 => L2_n_30, A3 => L2_n_134, B => L2_n_153, ZN => L2_n_158);
  L2_g7567 : OAI32D1BWP7T port map(A1 => L2_vgacontrol_vcount(9), A2 => L2_n_88, A3 => L2_n_134, B1 => L2_n_5, B2 => L2_n_137, ZN => L2_n_157);
  L2_g7568 : OAI32D1BWP7T port map(A1 => L2_vgacontrol_vcount(4), A2 => L2_n_521, A3 => L2_n_134, B1 => L2_n_6, B2 => L2_n_140, ZN => L2_n_156);
  L2_g7569 : MOAI22D0BWP7T port map(A1 => L2_n_127, A2 => L2_current_block_horizontal(3), B1 => L2_n_127, B2 => L2_current_block_horizontal(3), ZN => L2_n_155);
  L2_g7570 : ND2D1BWP7T port map(A1 => L2_n_141, A2 => L2_vgacontrol_vcount(6), ZN => L2_n_153);
  L2_g7571 : OAI21D0BWP7T port map(A1 => L2_n_132, A2 => L2_n_76, B => L2_vgacontrol_vcount(8), ZN => L2_n_152);
  L2_g7572 : OAI21D0BWP7T port map(A1 => L2_n_132, A2 => L2_n_26, B => L2_vgacontrol_vcount(1), ZN => L2_n_151);
  L2_g7573 : IND2D1BWP7T port map(A1 => L2_n_127, B1 => L2_current_block_horizontal(3), ZN => L2_n_154);
  L2_g7576 : AO21D0BWP7T port map(A1 => L2_n_125, A2 => L2_n_3, B => L2_n_144, Z => L2_n_150);
  L2_g7577 : OAI21D0BWP7T port map(A1 => L2_vgacontrol_vcount(4), A2 => L2_n_1, B => L2_n_140, ZN => L2_n_149);
  L2_g7578 : AO21D0BWP7T port map(A1 => L2_n_10, A2 => L2_n_2, B => L2_n_141, Z => L2_n_148);
  L2_g7579 : AOI21D0BWP7T port map(A1 => L2_n_130, A2 => L2_n_523, B => L2_n_1, ZN => L2_n_147);
  L2_g7580 : OAI32D1BWP7T port map(A1 => L2_vgacontrol_vcount(0), A2 => L2_n_121, A3 => L2_n_134, B1 => L2_n_4, B2 => L2_n_133, ZN => L2_n_146);
  L2_g7581 : MOAI22D0BWP7T port map(A1 => L2_n_123, A2 => L2_vgacontrol_hcount(9), B1 => L2_n_123, B2 => L2_vgacontrol_hcount(9), ZN => L2_n_145);
  L2_g7582 : NR4D0BWP7T port map(A1 => L2_n_134, A2 => L2_n_521, A3 => L2_n_6, A4 => L2_vgacontrol_vcount(5), ZN => L2_n_142);
  L2_g7583 : IOA21D1BWP7T port map(A1 => L2_n_125, A2 => L2_n_525, B => L2_n_133, ZN => L2_n_144);
  L2_g7584 : INR3D0BWP7T port map(A1 => L2_n_125, B1 => L2_n_525, B2 => L2_n_126, ZN => L2_n_143);
  L2_g7587 : OR4D1BWP7T port map(A1 => L2_vgacontrol_vcount(7), A2 => L2_n_10, A3 => L2_n_30, A4 => L2_n_134, Z => L2_n_139);
  L2_g7588 : OAI21D0BWP7T port map(A1 => L2_n_122, A2 => L2_n_524, B => L2_n_131, ZN => L2_n_138);
  L2_g7589 : AOI21D0BWP7T port map(A1 => L2_n_125, A2 => L2_n_88, B => L2_n_132, ZN => L2_n_137);
  L2_g7590 : MOAI22D0BWP7T port map(A1 => L2_n_118, A2 => L2_current_block_vertical(3), B1 => L2_n_118, B2 => L2_current_block_vertical(3), ZN => L2_n_136);
  L2_g7591 : IOA21D1BWP7T port map(A1 => L2_n_30, A2 => L2_n_2, B => L2_n_133, ZN => L2_n_141);
  L2_g7592 : AOI21D0BWP7T port map(A1 => L2_n_521, A2 => L2_n_2, B => L2_n_132, ZN => L2_n_140);
  L2_g7593 : IND2D1BWP7T port map(A1 => L2_n_118, B1 => L2_current_block_vertical(3), ZN => L2_n_135);
  L2_g7596 : OR2D1BWP7T port map(A1 => L2_n_126, A2 => L2_n_1, Z => L2_n_134);
  L2_g7597 : INVD1BWP7T port map(I => L2_n_133, ZN => L2_n_132);
  L2_g7598 : OAI21D0BWP7T port map(A1 => L2_n_122, A2 => L2_n_32, B => L2_n_12, ZN => L2_n_131);
  L2_g7599 : OAI31D0BWP7T port map(A1 => L2_n_97, A2 => L2_n_105, A3 => L2_n_120, B => calc_start_game_int, ZN => L2_n_130);
  L2_g7600 : MOAI22D0BWP7T port map(A1 => L2_n_111, A2 => L2_current_block_horizontal(2), B1 => L2_n_111, B2 => L2_current_block_horizontal(2), ZN => L2_n_129);
  L2_g7601 : MOAI22D0BWP7T port map(A1 => L2_n_112, A2 => L2_county(2), B1 => L2_n_112, B2 => L2_county(2), ZN => L2_n_128);
  L2_g7602 : ND2D1BWP7T port map(A1 => L2_n_126, A2 => L2_n_2, ZN => L2_n_133);
  L2_g7609 : MOAI22D0BWP7T port map(A1 => L2_n_104, A2 => L2_vgacontrol_hcount(8), B1 => L2_n_104, B2 => L2_vgacontrol_hcount(8), ZN => L2_n_124);
  L2_g7610 : IND2D1BWP7T port map(A1 => L2_n_111, B1 => L2_current_block_horizontal(2), ZN => L2_n_127);
  L2_g7611 : IND4D0BWP7T port map(A1 => L2_vgacontrol_hcount(7), B1 => L2_vgacontrol_hcount(4), B2 => L2_vgacontrol_hcount(6), B3 => L2_n_109, ZN => L2_n_126);
  L2_g7612 : NR2D1BWP7T port map(A1 => L2_n_121, A2 => L2_n_1, ZN => L2_n_125);
  L2_g7615 : IND2D1BWP7T port map(A1 => L2_n_104, B1 => L2_vgacontrol_hcount(8), ZN => L2_n_123);
  L2_g7618 : INVD0BWP7T port map(I => L2_n_120, ZN => L2_n_121);
  L2_g7619 : MOAI22D0BWP7T port map(A1 => L2_n_96, A2 => L2_current_block_vertical(2), B1 => L2_n_96, B2 => L2_current_block_vertical(2), ZN => L2_n_119);
  L2_g7620 : IND3D1BWP7T port map(A1 => L2_vgacontrol_hcount(7), B1 => L2_vgacontrol_hcount(6), B2 => L2_n_108, ZN => L2_n_122);
  L2_g7621 : ND4D0BWP7T port map(A1 => L2_n_103, A2 => L2_n_6, A3 => L2_n_4, A4 => L2_vgacontrol_vcount(2), ZN => L2_n_120);
  L2_g7627 : MOAI22D0BWP7T port map(A1 => L2_n_530, A2 => L2_calc_start_internal, B1 => L2_n_95, B2 => L2_n_100, ZN => L2_n_116);
  L2_g7628 : MOAI22D0BWP7T port map(A1 => L2_n_86, A2 => L2_current_block_horizontal(1), B1 => L2_n_86, B2 => L2_current_block_horizontal(1), ZN => L2_n_115);
  L2_g7629 : MOAI22D0BWP7T port map(A1 => L2_n_87, A2 => L2_in_go_y_pos(1), B1 => L2_n_87, B2 => L2_in_go_y_pos(1), ZN => L2_n_114);
  L2_g7630 : NR4D0BWP7T port map(A1 => L2_n_94, A2 => L2_n_4, A3 => L2_vgacontrol_vcount(4), A4 => L2_vgacontrol_vcount(2), ZN => L2_n_113);
  L2_g7631 : IND2D1BWP7T port map(A1 => L2_n_96, B1 => L2_current_block_vertical(2), ZN => L2_n_118);
  L2_g7632 : OA21D0BWP7T port map(A1 => L2_n_105, A2 => L2_n_31, B => L2_n_2, Z => L2_n_117);
  L2_g7633 : IND2D1BWP7T port map(A1 => L2_n_87, B1 => L2_in_go_y_pos(1), ZN => L2_n_112);
  L2_g7636 : IND2D1BWP7T port map(A1 => L2_n_86, B1 => L2_current_block_horizontal(1), ZN => L2_n_111);
  L2_g7637 : OAI22D0BWP7T port map(A1 => L2_n_91, A2 => L2_n_1, B1 => game_over_out_int, B2 => L2_n_42, ZN => L2_n_110);
  L2_g7638 : AN4D0BWP7T port map(A1 => L2_n_78, A2 => L2_vgacontrol_hcount(0), A3 => L2_vgacontrol_hcount(2), A4 => L2_vgacontrol_hcount(3), Z => L2_n_109);
  L2_g7639 : NR3D0BWP7T port map(A1 => L2_n_97, A2 => L2_n_22, A3 => L2_vgacontrol_hcount(3), ZN => L2_n_108);
  L2_g7640 : MOAI22D0BWP7T port map(A1 => L2_n_49, A2 => L2_vgacontrol_hcount(7), B1 => L2_n_49, B2 => L2_vgacontrol_hcount(7), ZN => L2_n_107);
  L2_g7641 : AO22D0BWP7T port map(A1 => L2_n_95, A2 => L2_n_39, B1 => L2_shift_L12_count_internal(1), B2 => L2_n_33, Z => L2_n_106);
  L2_g7642 : NR4D0BWP7T port map(A1 => L2_n_37, A2 => L2_n_5, A3 => L2_vgacontrol_vcount(8), A4 => L2_vgacontrol_vcount(7), ZN => L2_n_103);
  L2_g7643 : IND4D0BWP7T port map(A1 => L2_vgacontrol_hcount(6), B1 => L2_vgacontrol_hcount(3), B2 => L2_vgacontrol_hcount(7), B3 => L2_n_44, ZN => L2_n_105);
  L2_g7644 : IND2D1BWP7T port map(A1 => L2_n_49, B1 => L2_vgacontrol_hcount(7), ZN => L2_n_104);
  L2_g7647 : MOAI22D0BWP7T port map(A1 => L2_n_31, A2 => L2_vgacontrol_hcount(3), B1 => L2_n_31, B2 => L2_vgacontrol_hcount(3), ZN => L2_n_102);
  L2_g7648 : MOAI22D0BWP7T port map(A1 => L2_n_21, A2 => L2_current_block_vertical(1), B1 => L2_n_21, B2 => L2_current_block_vertical(1), ZN => L2_n_101);
  L2_g7649 : MOAI22D0BWP7T port map(A1 => L2_n_25, A2 => L2_shift_L12_count_internal(2), B1 => L2_n_25, B2 => L2_shift_L12_count_internal(2), ZN => L2_n_100);
  L2_g7650 : MOAI22D0BWP7T port map(A1 => L2_n_24, A2 => L2_vgacontrol_hcount(5), B1 => L2_n_24, B2 => L2_vgacontrol_hcount(5), ZN => L2_n_99);
  L2_g7651 : MOAI22D0BWP7T port map(A1 => L2_n_89, A2 => L2_n_533, B1 => L2_n_89, B2 => L2_screencontrol_go, ZN => L2_n_98);
  L2_g7671 : ND4D0BWP7T port map(A1 => L2_n_17, A2 => L2_n_5, A3 => L2_vgacontrol_vcount(7), A4 => L2_vgacontrol_vcount(8), ZN => L2_n_94);
  L2_g7672 : MOAI22D0BWP7T port map(A1 => L2_n_47, A2 => L2_county(0), B1 => L2_n_47, B2 => L2_county(0), ZN => L2_n_93);
  L2_g7673 : MOAI22D0BWP7T port map(A1 => L2_n_40, A2 => L2_current_block_horizontal(0), B1 => L2_n_40, B2 => L2_current_block_horizontal(0), ZN => L2_n_92);
  L2_g7674 : AOI211XD0BWP7T port map(A1 => L2_screencontrol_n_66, A2 => L2_n_16, B => L2_n_45, C => L2_in_st_go_sel, ZN => L2_n_91);
  L2_g7675 : MOAI22D0BWP7T port map(A1 => L2_n_14, A2 => L2_n_42, B1 => L2_n_43, B2 => L2_n_2, ZN => L2_n_90);
  L2_g7686 : ND3D0BWP7T port map(A1 => L2_vgacontrol_hcount(0), A2 => L2_vgacontrol_hcount(1), A3 => L2_vgacontrol_hcount(2), ZN => L2_n_97);
  L2_g7688 : IND2D1BWP7T port map(A1 => L2_n_21, B1 => L2_current_block_vertical(1), ZN => L2_n_96);
  L2_g7689 : CKAN2D1BWP7T port map(A1 => L2_n_79, A2 => L2_calc_start_internal, Z => L2_n_95);
  L2_g7690 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_x(1), B1 => L2_shift_pacman_pos_x_new(1), B2 => L2_n_29, Z => L2_n_85);
  L2_g7691 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_x(0), B1 => L2_shift_gr_pos_x_new(0), B2 => L2_n_28, Z => L2_n_84);
  L2_g7692 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_y(4), B1 => L2_shift_pacman_pos_y_new(4), B2 => L2_n_29, Z => L2_n_83);
  L2_g7693 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_y(3), B1 => L2_shift_pacman_pos_y_new(3), B2 => L2_n_29, Z => L2_n_82);
  L2_g7694 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_y(2), B1 => L2_shift_pacman_pos_y_new(2), B2 => L2_n_29, Z => L2_n_81);
  L2_g7695 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_y(1), B1 => L2_shift_pacman_pos_y_new(1), B2 => L2_n_29, Z => L2_n_80);
  L2_g7696 : AOI31D0BWP7T port map(A1 => L2_n_8, A2 => L2_n_7, A3 => L2_shift_L12_count_internal(2), B => L2_shift_shift_clock_reset, ZN => L2_n_79);
  L2_g7697 : NR3D0BWP7T port map(A1 => L2_n_22, A2 => L2_vgacontrol_hcount(5), A3 => L2_vgacontrol_hcount(1), ZN => L2_n_78);
  L2_g7698 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_x(0), B1 => L2_shift_pacman_pos_x_new(0), B2 => L2_n_29, Z => L2_n_77);
  L2_g7699 : AN2D0BWP7T port map(A1 => L2_n_48, A2 => L2_n_2, Z => L2_n_76);
  L2_g7700 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_x(2), B1 => L2_shift_pacman_pos_x_new(2), B2 => L2_n_29, Z => L2_n_75);
  L2_g7701 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_x(3), B1 => L2_shift_pacman_pos_x_new(3), B2 => L2_n_29, Z => L2_n_74);
  L2_g7702 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_x(4), B1 => L2_shift_pacman_pos_x_new(4), B2 => L2_n_29, Z => L2_n_73);
  L2_g7703 : AO22D0BWP7T port map(A1 => L2_n_27, A2 => L2_shift_pacman_pos_y(0), B1 => L2_shift_pacman_pos_y_new(0), B2 => L2_n_29, Z => L2_n_72);
  L2_g7704 : AOI31D0BWP7T port map(A1 => game_over_out_int, A2 => L2_n_11, A3 => L2_screencontrol_state(0), B => L2_n_533, ZN => L2_n_89);
  L2_g7705 : INR4D0BWP7T port map(A1 => L2_n_41, B1 => L2_en_dual_pixel_y_video, B2 => L2_en_dual_pixel_y_go, B3 => L2_en_dual_pixel_y_score, ZN => L2_n_71);
  L2_g7706 : IND2D1BWP7T port map(A1 => L2_n_48, B1 => L2_vgacontrol_vcount(8), ZN => L2_n_88);
  L2_g7707 : IND2D1BWP7T port map(A1 => L2_n_47, B1 => L2_county(0), ZN => L2_n_87);
  L2_g7708 : IND2D1BWP7T port map(A1 => L2_n_40, B1 => L2_current_block_horizontal(0), ZN => L2_n_86);
  L2_g7709 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_x(1), B1 => L2_shift_gr_pos_x_new(1), B2 => L2_n_28, Z => L2_n_70);
  L2_g7710 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_x(2), B1 => L2_shift_gr_pos_x_new(2), B2 => L2_n_28, Z => L2_n_69);
  L2_g7711 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_x(3), B1 => L2_shift_gr_pos_x_new(3), B2 => L2_n_28, Z => L2_n_68);
  L2_g7712 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_x(4), B1 => L2_shift_gr_pos_x_new(4), B2 => L2_n_28, Z => L2_n_67);
  L2_g7713 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_y(0), B1 => L2_shift_gr_pos_y_new(0), B2 => L2_n_28, Z => L2_n_66);
  L2_g7714 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_y(1), B1 => L2_shift_gr_pos_y_new(1), B2 => L2_n_28, Z => L2_n_65);
  L2_g7715 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_y(2), B1 => L2_shift_gr_pos_y_new(2), B2 => L2_n_28, Z => L2_n_64);
  L2_g7716 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_y(3), B1 => L2_shift_gr_pos_y_new(3), B2 => L2_n_28, Z => L2_n_63);
  L2_g7717 : AO22D0BWP7T port map(A1 => L2_n_19, A2 => L2_shift_gr_pos_y(4), B1 => L2_shift_gr_pos_y_new(4), B2 => L2_n_28, Z => L2_n_62);
  L2_g7718 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_x(0), B1 => L2_shift_gg_pos_x_new(0), B2 => L2_n_18, Z => L2_n_61);
  L2_g7719 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_x(1), B1 => L2_shift_gg_pos_x_new(1), B2 => L2_n_18, Z => L2_n_60);
  L2_g7720 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_x(2), B1 => L2_shift_gg_pos_x_new(2), B2 => L2_n_18, Z => L2_n_59);
  L2_g7721 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_x(3), B1 => L2_shift_gg_pos_x_new(3), B2 => L2_n_18, Z => L2_n_58);
  L2_g7722 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_x(4), B1 => L2_shift_gg_pos_x_new(4), B2 => L2_n_18, Z => L2_n_57);
  L2_g7723 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_y(0), B1 => L2_shift_gg_pos_y_new(0), B2 => L2_n_18, Z => L2_n_56);
  L2_g7724 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_y(1), B1 => L2_shift_gg_pos_y_new(1), B2 => L2_n_18, Z => L2_n_55);
  L2_g7725 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_y(2), B1 => L2_shift_gg_pos_y_new(2), B2 => L2_n_18, Z => L2_n_54);
  L2_g7726 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_y(3), B1 => L2_shift_gg_pos_y_new(3), B2 => L2_n_18, Z => L2_n_53);
  L2_g7727 : AO22D0BWP7T port map(A1 => L2_n_20, A2 => L2_shift_gg_pos_y(4), B1 => L2_shift_gg_pos_y_new(4), B2 => L2_n_18, Z => L2_n_52);
  L2_g7728 : MOAI22D0BWP7T port map(A1 => L2_n_23, A2 => L2_vgacontrol_hcount(6), B1 => L2_n_23, B2 => L2_vgacontrol_hcount(6), ZN => L2_n_51);
  L2_g7729 : INR3D0BWP7T port map(A1 => L2_screencontrol_n_58, B1 => L2_screencontrol_state(1), B2 => L2_screencontrol_state(0), ZN => L2_n_45);
  L2_g7730 : NR2XD0BWP7T port map(A1 => L2_n_32, A2 => L2_n_22, ZN => L2_n_44);
  L2_g7731 : OAI21D0BWP7T port map(A1 => L2_screencontrol_n_58, A2 => L2_n_15, B => L2_n_532, ZN => L2_n_43);
  L2_g7732 : NR3D0BWP7T port map(A1 => L2_reset_county_go, A2 => L2_reset_county_score, A3 => L2_reset_county_video, ZN => L2_n_50);
  L2_g7733 : IND2D1BWP7T port map(A1 => L2_n_23, B1 => L2_vgacontrol_hcount(6), ZN => L2_n_49);
  L2_g7734 : OR2D1BWP7T port map(A1 => L2_n_30, A2 => L2_n_522, Z => L2_n_48);
  L2_g7735 : NR3D0BWP7T port map(A1 => L2_en_county_go, A2 => L2_en_county_score, A3 => L2_en_county_video, ZN => L2_n_47);
  L2_g7736 : NR3D0BWP7T port map(A1 => L2_reset_current_block_horizontal_go, A2 => L2_reset_current_block_horizontal_score, A3 => L2_reset_current_block_horizontal_video, ZN => L2_n_46);
  L2_g7737 : OAI22D0BWP7T port map(A1 => L2_n_7, A2 => L2_shift_L12_count_internal(1), B1 => L2_n_8, B2 => L2_shift_L12_count_internal(0), ZN => L2_n_39);
  L2_g7738 : MOAI22D0BWP7T port map(A1 => L2_n_526, A2 => L2_vgacontrol_hcount(4), B1 => L2_n_526, B2 => L2_vgacontrol_hcount(4), ZN => L2_n_38);
  L2_g7739 : IND3D1BWP7T port map(A1 => L2_vgacontrol_vcount(1), B1 => L2_vgacontrol_vcount(3), B2 => L2_n_528, ZN => L2_n_37);
  L2_g7740 : CKXOR2D1BWP7T port map(A1 => L2_n_527, A2 => L2_vgacontrol_hcount(2), Z => L2_n_36);
  L2_g7741 : CKXOR2D1BWP7T port map(A1 => L2_en_current_block_vertical, A2 => L2_current_block_vertical(0), Z => L2_n_35);
  L2_g7742 : MOAI22D0BWP7T port map(A1 => L2_n_9, A2 => L2_vgacontrol_hcount(1), B1 => L2_n_9, B2 => L2_vgacontrol_hcount(1), ZN => L2_n_34);
  L2_g7743 : ND3D0BWP7T port map(A1 => L2_n_11, A2 => L2_screencontrol_state(0), A3 => L2_n_2, ZN => L2_n_42);
  L2_g7744 : NR3D0BWP7T port map(A1 => L2_reset_dual_pixel_y_go, A2 => L2_reset_dual_pixel_y_score, A3 => L2_reset_dual_pixel_y_video, ZN => L2_n_41);
  L2_g7745 : NR3D0BWP7T port map(A1 => L2_en_current_block_horizontal_go, A2 => L2_en_current_block_horizontal_score, A3 => L2_en_current_block_horizontal_video, ZN => L2_n_40);
  L2_g7746 : NR2XD0BWP7T port map(A1 => L2_vgacontrol_vcount(0), A2 => L2_n_1, ZN => L2_n_26);
  L2_g7747 : NR2D1BWP7T port map(A1 => L2_shift_shift_clock_reset, A2 => L2_calc_start_internal, ZN => L2_n_33);
  L2_g7748 : OR2D1BWP7T port map(A1 => L2_vgacontrol_hcount(5), A2 => L2_vgacontrol_hcount(4), Z => L2_n_32);
  L2_g7749 : ND2D1BWP7T port map(A1 => L2_n_527, A2 => L2_vgacontrol_hcount(2), ZN => L2_n_31);
  L2_g7750 : IND2D1BWP7T port map(A1 => L2_n_521, B1 => L2_n_529, ZN => L2_n_30);
  L2_g7751 : INR2XD0BWP7T port map(A1 => L2_shift_pacman_pos_load, B1 => L2_shift_pacman_pos_reset, ZN => L2_n_29);
  L2_g7752 : INR2XD0BWP7T port map(A1 => L2_shift_gr_pos_load, B1 => L2_shift_gr_pos_reset, ZN => L2_n_28);
  L2_g7753 : NR2XD0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => L2_shift_pacman_pos_reset, ZN => L2_n_27);
  L2_g7754 : INR2XD0BWP7T port map(A1 => L2_vgacontrol_vcount(3), B1 => L2_n_552, ZN => L2_n_17);
  L2_g7755 : CKND2D1BWP7T port map(A1 => L2_shift_L12_count_internal(0), A2 => L2_shift_L12_count_internal(1), ZN => L2_n_25);
  L2_g7756 : IND2D1BWP7T port map(A1 => L2_n_526, B1 => L2_vgacontrol_hcount(4), ZN => L2_n_24);
  L2_g7757 : OR2D1BWP7T port map(A1 => L2_n_526, A2 => L2_n_524, Z => L2_n_23);
  L2_g7758 : IND2D1BWP7T port map(A1 => L2_vgacontrol_hcount(9), B1 => L2_vgacontrol_hcount(8), ZN => L2_n_22);
  L2_g7759 : ND2D1BWP7T port map(A1 => L2_en_current_block_vertical, A2 => L2_current_block_vertical(0), ZN => L2_n_21);
  L2_g7760 : NR2XD0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => L2_shift_gg_pos_reset, ZN => L2_n_20);
  L2_g7761 : NR2XD0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => L2_shift_gr_pos_reset, ZN => L2_n_19);
  L2_g7762 : INR2XD0BWP7T port map(A1 => L2_shift_gg_pos_load, B1 => L2_shift_gg_pos_reset, ZN => L2_n_18);
  L2_g7806 : CKND1BWP7T port map(I => L2_n_532, ZN => L2_n_16);
  L2_g7807 : INVD1BWP7T port map(I => L2_in_st_go_sel, ZN => L2_n_15);
  L2_g7808 : INVD0BWP7T port map(I => game_over_out_int, ZN => L2_n_14);
  L2_g7825 : INVD1BWP7T port map(I => L2_reset_current_block_vertical, ZN => L2_n_13);
  L2_screencontrol_state_reg_1 : DFD1BWP7T port map(CP => clk, D => L2_n_90, Q => L2_screencontrol_state(1), QN => L2_n_11);
  L2_shift_L12_count_internal_reg_0 : DFXD1BWP7T port map(CP => clk, DA => L2_n_33, DB => L2_n_95, SA => L2_shift_L12_count_internal(0), Q => L2_shift_L12_count_internal(0), QN => L2_n_7);
  L2_shift_L12_count_internal_reg_1 : DFD1BWP7T port map(CP => clk, D => L2_n_106, Q => L2_shift_L12_count_internal(1), QN => L2_n_8);
  L2_vgacontrol_hcount_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => L2_n_9, D => L2_n_117, Q => L2_vgacontrol_hcount(0), QN => L2_n_9);
  L2_vgacontrol_in_h_sync_reg : DFKCND0BWP7T port map(CP => clk, CN => L2_n_2, D => L2_n_138, Q => L2_n_12, QN => L2_n_0);
  L2_vgacontrol_vcount_reg_0 : DFD1BWP7T port map(CP => clk, D => L2_n_146, Q => L2_vgacontrol_vcount(0), QN => L2_n_4);
  L2_vgacontrol_vcount_reg_2 : DFXD1BWP7T port map(CP => clk, DA => L2_n_144, DB => L2_n_143, SA => L2_vgacontrol_vcount(2), Q => L2_vgacontrol_vcount(2), QN => L2_n_3);
  L2_vgacontrol_vcount_reg_4 : DFD1BWP7T port map(CP => clk, D => L2_n_156, Q => L2_vgacontrol_vcount(4), QN => L2_n_6);
  L2_vgacontrol_vcount_reg_6 : DFD1BWP7T port map(CP => clk, D => L2_n_158, Q => L2_vgacontrol_vcount(6), QN => L2_n_10);
  L2_vgacontrol_vcount_reg_9 : DFD1BWP7T port map(CP => clk, D => L2_n_157, Q => L2_vgacontrol_vcount(9), QN => L2_n_5);
  L2_drc_bufs7851 : INVD1BWP7T port map(I => L2_n_2, ZN => L2_n_1);
  L2_drc_bufs7852 : INVD0BWP7T port map(I => reset, ZN => L2_n_2);
  L2_drc_bufs7855 : INVD4BWP7T port map(I => L2_n_0, ZN => h_sync);
  L2_drc_bufs7858 : BUFFD4BWP7T port map(I => L2_n_167, Z => v_sync);
  L2_cnt_in_county_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => L2_n_50, D => L2_n_128, Q => L2_county(2), QN => L2_n_230);
  L2_cnt_in_county_reg_1 : DFKCND1BWP7T port map(CP => clk, CN => L2_n_50, D => L2_n_114, Q => L2_in_go_y_pos(1), QN => L2_n_229);
  L2_cnt_in_county_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => L2_n_93, D => L2_n_50, Q => L2_county(0), QN => L2_n_226);
  L2_shift_L31_shift_sync_gg_reg : DFQD0BWP7T port map(CP => clk, D => L2_shift_L31_n_9, Q => L2_shift_shift_pulse_gg);
  L2_shift_L31_g174 : INR4D0BWP7T port map(A1 => L2_calc_start_internal, B1 => L2_shift_L31_count_internal(0), B2 => L2_shift_L31_n_8, B3 => L2_shift_shift_clock_reset_gg, ZN => L2_shift_L31_n_9);
  L2_shift_L31_g175 : IND2D1BWP7T port map(A1 => L2_shift_L31_count_internal(1), B1 => L2_shift_L31_count_internal(2), ZN => L2_shift_L31_n_8);
  L2_shift_L31_count_internal_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L31_n_7, Q => L2_shift_L31_count_internal(2));
  L2_shift_L31_count_internal_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L31_n_6, Q => L2_shift_L31_count_internal(1));
  L2_shift_L31_g244 : AO22D0BWP7T port map(A1 => L2_shift_L31_n_3, A2 => L2_shift_L31_n_4, B1 => L2_shift_L31_count_internal(2), B2 => L2_shift_L31_n_1, Z => L2_shift_L31_n_7);
  L2_shift_L31_g246 : AO22D0BWP7T port map(A1 => L2_shift_L31_n_3, A2 => L2_shift_L31_n_2, B1 => L2_shift_L31_count_internal(1), B2 => L2_shift_L31_n_1, Z => L2_shift_L31_n_6);
  L2_shift_L31_g247 : AO22D0BWP7T port map(A1 => L2_shift_L31_n_3, A2 => L2_shift_L31_n_10, B1 => L2_shift_L31_count_internal(0), B2 => L2_shift_L31_n_1, Z => L2_shift_L31_n_5);
  L2_shift_L31_g248 : MOAI22D0BWP7T port map(A1 => L2_shift_L31_n_0, A2 => L2_shift_L31_count_internal(2), B1 => L2_shift_L31_n_0, B2 => L2_shift_L31_count_internal(2), ZN => L2_shift_L31_n_4);
  L2_shift_L31_g249 : NR3D0BWP7T port map(A1 => L2_shift_L31_n_9, A2 => L2_shift_L31_n_1, A3 => L2_shift_shift_clock_reset_gg, ZN => L2_shift_L31_n_3);
  L2_shift_L31_g250 : MOAI22D0BWP7T port map(A1 => L2_shift_L31_n_10, A2 => L2_shift_L31_count_internal(1), B1 => L2_shift_L31_n_10, B2 => L2_shift_L31_count_internal(1), ZN => L2_shift_L31_n_2);
  L2_shift_L31_g251 : NR2XD0BWP7T port map(A1 => L2_shift_shift_clock_reset_gg, A2 => L2_calc_start_internal, ZN => L2_shift_L31_n_1);
  L2_shift_L31_g252 : ND2D1BWP7T port map(A1 => L2_shift_L31_count_internal(1), A2 => L2_shift_L31_count_internal(0), ZN => L2_shift_L31_n_0);
  L2_shift_L31_count_internal_reg_0 : DFD1BWP7T port map(CP => clk, D => L2_shift_L31_n_5, Q => L2_shift_L31_count_internal(0), QN => L2_shift_L31_n_10);
  L2_shift_L33_g12867 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_272, A2 => L2_county(0), B => L2_shift_L33_n_278, ZN => L2_shift_y_pos_out_shift_gg(0));
  L2_shift_L33_g12868 : OR4D1BWP7T port map(A1 => L2_shift_L33_n_264, A2 => L2_shift_L33_n_268, A3 => L2_shift_L33_n_267, A4 => L2_shift_L33_n_276, Z => L2_shift_y_pos_out_shift_gg(2));
  L2_shift_L33_g12869 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_175, A2 => L2_shift_L33_n_269, B => L2_shift_L33_n_277, C => L2_shift_L33_n_270, ZN => L2_shift_y_pos_out_shift_gg(1));
  L2_shift_L33_g12870 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_275, A2 => L2_shift_L33_n_266, B => L2_county(0), ZN => L2_shift_L33_n_278);
  L2_shift_L33_g12871 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_275, A2 => L2_in_go_y_pos(1), B1 => L2_shift_L33_n_265, B2 => L2_shift_L33_n_175, ZN => L2_shift_L33_n_277);
  L2_shift_L33_g12872 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_274, A2 => L2_shift_L33_n_52, B1 => L2_shift_L33_n_328, B2 => L2_shift_L33_n_302, ZN => L2_shift_L33_n_276);
  L2_shift_L33_g12873 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_283, B1 => L2_shift_L33_n_274, ZN => L2_shift_L33_n_275);
  L2_shift_L33_g12874 : IIND4D0BWP7T port map(A1 => L2_shift_L33_n_265, A2 => L2_shift_L33_n_286, B1 => L2_shift_L33_n_273, B2 => L2_shift_L33_n_252, ZN => L2_shift_L33_n_274);
  L2_shift_L33_g12875 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_266, A2 => L2_shift_L33_n_280, A3 => L2_shift_L33_n_283, A4 => L2_shift_L33_n_282, ZN => L2_shift_L33_n_273);
  L2_shift_L33_g12876 : CKAN2D1BWP7T port map(A1 => cell_type_int(2), A2 => L2_shift_L33_n_271, Z => L2_shift_cell_state_out_shift_gg(2));
  L2_shift_L33_g12877 : IND2D1BWP7T port map(A1 => cell_type_int(1), B1 => L2_shift_L33_n_271, ZN => L2_shift_cell_state_out_shift_gg(1));
  L2_shift_L33_g12878 : IND2D1BWP7T port map(A1 => cell_type_int(0), B1 => L2_shift_L33_n_271, ZN => L2_shift_cell_state_out_shift_gg(0));
  L2_shift_L33_g12879 : INR2XD0BWP7T port map(A1 => L2_shift_L33_n_269, B1 => L2_shift_L33_n_265, ZN => L2_shift_L33_n_272);
  L2_shift_L33_g12880 : AO21D0BWP7T port map(A1 => L2_shift_L33_n_258, A2 => L2_shift_L33_n_254, B => L2_in_go_y_pos(1), Z => L2_shift_L33_n_270);
  L2_shift_L33_g12881 : IND4D0BWP7T port map(A1 => L2_shift_L33_n_288, B1 => L2_shift_L33_n_247, B2 => L2_shift_L33_n_243, B3 => L2_shift_L33_n_250, ZN => L2_shift_L33_n_271);
  L2_shift_L33_g12882 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_258, A2 => L2_shift_L33_n_174, B => L2_shift_L33_n_263, ZN => L2_shift_L33_n_268);
  L2_shift_L33_g12883 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_261, A2 => L2_shift_L33_n_201, B1 => L2_shift_L33_n_259, B2 => L2_shift_L33_n_200, ZN => L2_shift_L33_n_267);
  L2_shift_L33_g12884 : INR3D0BWP7T port map(A1 => L2_shift_L33_n_252, B1 => L2_shift_L33_n_282, B2 => L2_shift_L33_n_262, ZN => L2_shift_L33_n_269);
  L2_shift_L33_g12885 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_260, A2 => L2_shift_L33_n_254, ZN => L2_shift_L33_n_266);
  L2_shift_L33_g12886 : OR2D1BWP7T port map(A1 => L2_shift_L33_n_259, A2 => L2_shift_L33_n_255, Z => L2_shift_L33_n_265);
  L2_shift_L33_g12887 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_256, A2 => L2_shift_L33_n_200, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_309, ZN => L2_shift_L33_n_264);
  L2_shift_L33_g12888 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_251, A2 => L2_shift_L33_n_201, B1 => L2_shift_L33_n_253, B2 => L2_shift_L33_n_174, ZN => L2_shift_L33_n_263);
  L2_shift_L33_g12889 : INVD1BWP7T port map(I => L2_shift_L33_n_261, ZN => L2_shift_L33_n_262);
  L2_shift_L33_g12890 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_285, A2 => L2_shift_L33_n_281, ZN => L2_shift_L33_n_260);
  L2_shift_L33_g12891 : IAO21D0BWP7T port map(A1 => L2_shift_L33_n_241, A2 => L2_shift_L33_n_297, B => L2_shift_L33_n_286, ZN => L2_shift_L33_n_261);
  L2_shift_L33_g12892 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_235, A2 => L2_shift_L33_n_295, B => L2_shift_L33_n_257, ZN => L2_shift_L33_n_259);
  L2_shift_L33_g12893 : AOI21D0BWP7T port map(A1 => L2_shift_L33_n_245, A2 => L2_shift_L33_n_53, B => L2_shift_L33_n_285, ZN => L2_shift_L33_n_258);
  L2_shift_L33_g12895 : INVD0BWP7T port map(I => L2_shift_L33_n_255, ZN => L2_shift_L33_n_256);
  L2_shift_L33_g12896 : INVD0BWP7T port map(I => L2_shift_L33_n_254, ZN => L2_shift_L33_n_253);
  L2_shift_L33_g12897 : INVD0BWP7T port map(I => L2_shift_L33_n_252, ZN => L2_shift_L33_n_251);
  L2_shift_L33_g12898 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_236, A2 => L2_shift_L33_n_295, ZN => L2_shift_L33_n_257);
  L2_shift_L33_g12899 : INR2XD0BWP7T port map(A1 => L2_shift_L33_n_293, B1 => L2_shift_L33_n_244, ZN => L2_shift_L33_n_255);
  L2_shift_L33_g12900 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_238, A2 => L2_shift_L33_n_294, ZN => L2_shift_L33_n_254);
  L2_shift_L33_g12901 : CKAN2D1BWP7T port map(A1 => L2_shift_L33_n_246, A2 => L2_shift_L33_n_297, Z => L2_shift_L33_n_286);
  L2_shift_L33_g12902 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_249, B1 => L2_shift_L33_n_279, ZN => L2_shift_L33_n_252);
  L2_shift_L33_g12903 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_289, A2 => L2_shift_L33_n_225, B1 => L2_shift_L33_n_290, B2 => L2_shift_L33_n_199, ZN => L2_shift_L33_n_250);
  L2_shift_L33_g12904 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_239, A2 => L2_shift_L33_n_294, ZN => L2_shift_L33_n_281);
  L2_shift_L33_g12905 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_240, A2 => L2_shift_L33_n_293, ZN => L2_shift_L33_n_280);
  L2_shift_L33_g12906 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_242, A2 => L2_shift_L33_n_53, ZN => L2_shift_L33_n_285);
  L2_shift_L33_g12907 : CKAN2D1BWP7T port map(A1 => L2_shift_L33_n_248, A2 => L2_county(2), Z => L2_shift_L33_n_283);
  L2_shift_L33_g12908 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_237, A2 => L2_shift_L33_n_279, ZN => L2_shift_L33_n_282);
  L2_shift_L33_g12909 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_328, A2 => L2_shift_L33_n_303, B1 => L2_shift_L33_n_227, B2 => L2_shift_L33_n_179, ZN => L2_shift_L33_n_249);
  L2_shift_L33_g12910 : AO22D0BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_309, B1 => L2_shift_L33_n_302, B2 => L2_shift_L33_n_298, Z => L2_shift_L33_n_248);
  L2_shift_L33_g12911 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_202, A2 => L2_shift_L33_n_320, B => L2_shift_L33_n_395, ZN => L2_shift_L33_n_247);
  L2_shift_L33_g12912 : AO22D0BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_312, B1 => L2_shift_L33_n_299, B2 => L2_shift_L33_n_298, Z => L2_shift_L33_n_246);
  L2_shift_L33_g12913 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_228, A2 => L2_shift_L33_n_184, B1 => L2_shift_L33_n_328, B2 => L2_shift_L33_n_300, ZN => L2_shift_L33_n_245);
  L2_shift_L33_g12914 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_328, A2 => L2_shift_L33_n_305, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_306, ZN => L2_shift_L33_n_244);
  L2_shift_L33_g12915 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_307, A2 => L2_shift_L33_n_218, B => L2_shift_L33_n_233, C => L2_shift_L33_n_219, ZN => L2_shift_L33_n_243);
  L2_shift_L33_g12916 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_311, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_300, ZN => L2_shift_L33_n_242);
  L2_shift_L33_g12917 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_328, A2 => L2_shift_L33_n_299, B1 => L2_shift_L33_n_227, B2 => L2_shift_L33_n_178, ZN => L2_shift_L33_n_241);
  L2_shift_L33_g12918 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_306, B1 => L2_shift_L33_n_227, B2 => L2_shift_L33_n_176, ZN => L2_shift_L33_n_240);
  L2_shift_L33_g12919 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_307, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_304, ZN => L2_shift_L33_n_239);
  L2_shift_L33_g12920 : AO22D0BWP7T port map(A1 => L2_shift_L33_n_328, A2 => L2_shift_L33_n_304, B1 => L2_shift_L33_n_307, B2 => L2_shift_L33_n_298, Z => L2_shift_L33_n_238);
  L2_shift_L33_g12921 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_308, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_303, ZN => L2_shift_L33_n_237);
  L2_shift_L33_g12922 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_228, A2 => L2_shift_L33_n_170, B1 => L2_shift_L33_n_393, B2 => L2_shift_L33_n_310, ZN => L2_shift_L33_n_236);
  L2_shift_L33_g12923 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_328, A2 => L2_shift_L33_n_301, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_310, ZN => L2_shift_L33_n_235);
  L2_shift_L33_g12925 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_298, ZN => L2_shift_L33_n_290);
  L2_shift_L33_g12926 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_328, A2 => L2_shift_L33_n_298, ZN => L2_shift_L33_n_289);
  L2_shift_L33_g12927 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_217, A2 => L2_shift_L33_n_231, A3 => L2_shift_L33_n_197, A4 => L2_shift_L33_n_209, ZN => L2_shift_L33_n_287);
  L2_shift_L33_g12928 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_216, A2 => L2_shift_L33_n_230, A3 => L2_shift_L33_n_198, A4 => L2_shift_L33_n_210, ZN => L2_shift_L33_n_328);
  L2_shift_L33_g12929 : INVD0BWP7T port map(I => L2_shift_L33_n_393, ZN => L2_shift_L33_n_233);
  L2_shift_L33_g12930 : INR4D0BWP7T port map(A1 => L2_shift_L33_n_197, B1 => L2_shift_L33_n_221, B2 => L2_shift_L33_n_232, B3 => L2_shift_L33_n_217, ZN => L2_shift_L33_n_394);
  L2_shift_L33_g12931 : INR4D0BWP7T port map(A1 => L2_shift_L33_n_198, B1 => L2_shift_L33_n_223, B2 => L2_shift_L33_n_229, B3 => L2_shift_L33_n_216, ZN => L2_shift_L33_n_393);
  L2_shift_L33_g12932 : OAI221D0BWP7T port map(A1 => L2_shift_L33_n_169, A2 => L2_shift_L33_n_207, B1 => L2_shift_L33_n_191, B2 => xcoordinates_int(2), C => L2_shift_L33_n_226, ZN => L2_shift_L33_n_232);
  L2_shift_L33_g12933 : OAI221D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L33_n_211, B1 => L2_shift_L33_n_208, B2 => L2_shift_L33_n_169, C => L2_shift_L33_n_222, ZN => L2_shift_L33_n_231);
  L2_shift_L33_g12934 : OAI221D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_L33_n_212, B1 => L2_shift_L33_n_204, B2 => L2_shift_L33_n_168, C => L2_shift_L33_n_220, ZN => L2_shift_L33_n_230);
  L2_shift_L33_g12935 : OAI221D0BWP7T port map(A1 => L2_shift_L33_n_168, A2 => L2_shift_L33_n_206, B1 => L2_shift_L33_n_192, B2 => ycoordinates_int(2), C => L2_shift_L33_n_224, ZN => L2_shift_L33_n_229);
  L2_shift_L33_g12936 : INVD0BWP7T port map(I => L2_shift_L33_n_228, ZN => L2_shift_L33_n_227);
  L2_shift_L33_g12937 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_169, A2 => L2_shift_L33_n_207, B1 => xcoordinates_int(2), B2 => L2_shift_L33_n_191, ZN => L2_shift_L33_n_226);
  L2_shift_L33_g12938 : OR4D1BWP7T port map(A1 => L2_shift_L33_n_299, A2 => L2_shift_L33_n_304, A3 => L2_shift_L33_n_302, A4 => L2_shift_L33_n_213, Z => L2_shift_L33_n_225);
  L2_shift_L33_g12939 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_168, A2 => L2_shift_L33_n_206, B1 => ycoordinates_int(2), B2 => L2_shift_L33_n_192, ZN => L2_shift_L33_n_224);
  L2_shift_L33_g12940 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_150, ZN => L2_shift_L33_n_228);
  L2_shift_L33_g12941 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_L33_n_215, B1 => ycoordinates_int(3), B2 => L2_shift_L33_n_215, ZN => L2_shift_L33_n_223);
  L2_shift_L33_g12942 : AOI22D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L33_n_211, B1 => L2_shift_L33_n_169, B2 => L2_shift_L33_n_208, ZN => L2_shift_L33_n_222);
  L2_shift_L33_g12943 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L33_n_214, B1 => xcoordinates_int(3), B2 => L2_shift_L33_n_214, ZN => L2_shift_L33_n_221);
  L2_shift_L33_g12944 : AOI22D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_L33_n_212, B1 => L2_shift_L33_n_168, B2 => L2_shift_L33_n_204, ZN => L2_shift_L33_n_220);
  L2_shift_L33_g12945 : INVD0BWP7T port map(I => L2_shift_L33_n_298, ZN => L2_shift_L33_n_219);
  L2_shift_L33_g12946 : AN4D1BWP7T port map(A1 => L2_shift_L33_n_203, A2 => L2_shift_L33_n_205, A3 => L2_shift_L33_n_168, A4 => L2_shift_L33_n_169, Z => L2_shift_L33_n_298);
  L2_shift_L33_g12947 : OR4D1BWP7T port map(A1 => L2_shift_L33_n_306, A2 => L2_shift_L33_n_309, A3 => L2_shift_L33_n_196, A4 => L2_shift_L33_n_310, Z => L2_shift_L33_n_218);
  L2_shift_L33_g12948 : ND3D0BWP7T port map(A1 => L2_shift_L33_n_203, A2 => L2_shift_L33_n_172, A3 => L2_shift_L33_n_168, ZN => L2_shift_L33_n_217);
  L2_shift_L33_g12949 : ND3D0BWP7T port map(A1 => L2_shift_L33_n_205, A2 => L2_shift_L33_n_173, A3 => L2_shift_L33_n_169, ZN => L2_shift_L33_n_216);
  L2_shift_L33_g12950 : AO211D0BWP7T port map(A1 => L2_shift_L33_n_195, A2 => L2_shift_L33_n_150, B => L2_shift_L33_n_300, C => L2_shift_L33_n_303, Z => L2_shift_L33_n_213);
  L2_shift_L33_g12951 : AOI21D0BWP7T port map(A1 => L2_shift_L33_n_187, A2 => L2_shift_gg_pos_y(3), B => L2_shift_L33_n_206, ZN => L2_shift_L33_n_215);
  L2_shift_L33_g12952 : AOI21D0BWP7T port map(A1 => L2_shift_L33_n_188, A2 => L2_shift_gg_pos_x(3), B => L2_shift_L33_n_207, ZN => L2_shift_L33_n_214);
  L2_shift_L33_g12953 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(2), A2 => L2_shift_L33_n_194, B1 => ycoordinates_int(2), B2 => L2_shift_L33_n_194, ZN => L2_shift_L33_n_210);
  L2_shift_L33_g12954 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(2), A2 => L2_shift_L33_n_193, B1 => xcoordinates_int(2), B2 => L2_shift_L33_n_193, ZN => L2_shift_L33_n_209);
  L2_shift_L33_g12955 : MAOI22D0BWP7T port map(A1 => L2_shift_L33_n_186, A2 => L2_shift_gg_pos_y(3), B1 => L2_shift_L33_n_186, B2 => L2_shift_gg_pos_y(3), ZN => L2_shift_L33_n_212);
  L2_shift_L33_g12956 : MAOI22D0BWP7T port map(A1 => L2_shift_L33_n_189, A2 => L2_shift_gg_pos_x(3), B1 => L2_shift_L33_n_189, B2 => L2_shift_gg_pos_x(3), ZN => L2_shift_L33_n_211);
  L2_shift_L33_g12957 : INR2D1BWP7T port map(A1 => L2_shift_gg_pos_x(3), B1 => L2_shift_L33_n_189, ZN => L2_shift_L33_n_208);
  L2_shift_L33_g12958 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_188, A2 => L2_shift_gg_pos_x(3), ZN => L2_shift_L33_n_207);
  L2_shift_L33_g12959 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_187, A2 => L2_shift_gg_pos_y(3), ZN => L2_shift_L33_n_206);
  L2_shift_L33_g12960 : OAI222D0BWP7T port map(A1 => L2_shift_L33_n_185, A2 => L2_shift_L33_n_150, B1 => L2_shift_L33_state(4), B2 => L2_shift_L33_n_180, C1 => L2_shift_L33_n_152, C2 => L2_shift_L33_n_156, ZN => L2_shift_L33_n_202);
  L2_shift_L33_g12961 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_172, A2 => L2_shift_L33_n_167, A3 => L2_shift_L33_n_143, A4 => L2_shift_L33_n_165, ZN => L2_shift_L33_n_205);
  L2_shift_L33_g12962 : INR2D1BWP7T port map(A1 => L2_shift_gg_pos_y(3), B1 => L2_shift_L33_n_186, ZN => L2_shift_L33_n_204);
  L2_shift_L33_g12963 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_171, A2 => L2_shift_L33_n_173, A3 => L2_shift_L33_n_166, A4 => L2_shift_L33_n_142, ZN => L2_shift_L33_n_203);
  L2_shift_L33_g12964 : OAI222D0BWP7T port map(A1 => L2_shift_L33_n_177, A2 => L2_shift_L33_n_152, B1 => L2_shift_L33_n_151, B2 => L2_shift_L33_n_156, C1 => L2_shift_L33_state(4), C2 => L2_shift_L33_n_160, ZN => L2_shift_L33_n_199);
  L2_shift_L33_g12965 : OA211D0BWP7T port map(A1 => L2_shift_L33_n_144, A2 => L2_shift_L33_n_52, B => L2_shift_L33_n_297, C => L2_shift_L33_n_294, Z => L2_shift_L33_n_201);
  L2_shift_L33_g12966 : OAI211D1BWP7T port map(A1 => L2_county(0), A2 => L2_county(2), B => L2_shift_L33_n_293, C => L2_shift_L33_n_296, ZN => L2_shift_L33_n_200);
  L2_shift_L33_g12967 : OAI21D0BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(0), B => L2_county(2), ZN => L2_shift_L33_n_279);
  L2_shift_L33_g12968 : AO21D0BWP7T port map(A1 => L2_shift_L33_n_150, A2 => L2_shift_L33_n_155, B => L2_shift_L33_n_308, Z => L2_shift_L33_n_196);
  L2_shift_L33_g12969 : MAOI22D0BWP7T port map(A1 => L2_shift_L33_n_171, A2 => L2_shift_gg_pos_y(0), B1 => L2_shift_L33_n_171, B2 => L2_shift_gg_pos_y(0), ZN => L2_shift_L33_n_198);
  L2_shift_L33_g12970 : MAOI22D0BWP7T port map(A1 => xcoordinates_int(1), A2 => L2_shift_L33_n_190, B1 => xcoordinates_int(1), B2 => L2_shift_L33_n_190, ZN => L2_shift_L33_n_197);
  L2_shift_L33_g12971 : AO21D0BWP7T port map(A1 => L2_shift_L33_n_181, A2 => L2_shift_L33_n_145, B => L2_shift_L33_n_387, Z => L2_shift_L33_n_288);
  L2_shift_L33_g12972 : IOA21D1BWP7T port map(A1 => L2_county(0), A2 => L2_in_go_y_pos(1), B => L2_shift_L33_n_52, ZN => L2_shift_L33_n_295);
  L2_shift_L33_g12973 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_183, A2 => L2_shift_L33_n_151, ZN => L2_shift_L33_n_318);
  L2_shift_L33_g12974 : INR2D1BWP7T port map(A1 => L2_shift_L33_state(1), B1 => L2_shift_L33_n_185, ZN => L2_shift_L33_n_321);
  L2_shift_L33_g12975 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_184, A2 => L2_shift_L33_n_152, ZN => L2_shift_L33_n_325);
  L2_shift_L33_g12976 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_183, A2 => L2_shift_L33_n_152, ZN => L2_shift_L33_n_316);
  L2_shift_L33_g12977 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_184, A2 => L2_shift_L33_n_151, ZN => L2_shift_L33_n_313);
  L2_shift_L33_g12978 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_178, B1 => L2_shift_L33_n_152, ZN => L2_shift_L33_n_326);
  L2_shift_L33_g12979 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_170, A2 => L2_shift_L33_n_177, ZN => L2_shift_L33_n_195);
  L2_shift_L33_g12980 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_180, A2 => L2_shift_L33_n_151, ZN => L2_shift_L33_n_324);
  L2_shift_L33_g12981 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_178, B1 => L2_shift_L33_n_151, ZN => L2_shift_L33_n_314);
  L2_shift_L33_g12982 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_180, A2 => L2_shift_L33_n_152, ZN => L2_shift_L33_n_322);
  L2_shift_L33_g12983 : CKAN2D1BWP7T port map(A1 => L2_shift_L33_n_178, A2 => L2_shift_L33_n_150, Z => L2_shift_L33_n_312);
  L2_shift_L33_g12984 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_184, A2 => L2_shift_L33_n_149, ZN => L2_shift_L33_n_311);
  L2_shift_L33_g12985 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_180, A2 => L2_shift_L33_n_149, ZN => L2_shift_L33_n_308);
  L2_shift_L33_g12986 : AN2D1BWP7T port map(A1 => L2_shift_L33_n_182, A2 => L2_shift_L33_n_150, Z => L2_shift_L33_n_302);
  L2_shift_L33_g12987 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_177, A2 => L2_shift_L33_n_154, ZN => L2_shift_L33_n_303);
  L2_shift_L33_g12988 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_183, A2 => L2_shift_L33_n_154, ZN => L2_shift_L33_n_300);
  L2_shift_L33_g12989 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_185, A2 => L2_shift_L33_n_145, ZN => L2_shift_L33_n_307);
  L2_shift_L33_g12990 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_181, B1 => L2_shift_L33_n_151, ZN => L2_shift_gg_pos_reset);
  L2_shift_L33_g12991 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_170, A2 => L2_shift_L33_n_151, ZN => L2_shift_L33_n_317);
  L2_shift_L33_g12992 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_170, A2 => L2_shift_L33_n_152, ZN => L2_shift_L33_n_315);
  L2_shift_L33_g12993 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_181, B1 => L2_shift_L33_n_152, ZN => L2_shift_L33_n_327);
  L2_shift_L33_g12994 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_185, A2 => L2_shift_L33_n_151, ZN => L2_shift_L33_n_323);
  L2_shift_L33_g12995 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_177, A2 => L2_shift_L33_n_151, ZN => L2_shift_L33_n_387);
  L2_shift_L33_g12996 : MAOI22D0BWP7T port map(A1 => L2_shift_L33_n_157, A2 => L2_shift_gg_pos_y(2), B1 => L2_shift_L33_n_157, B2 => L2_shift_gg_pos_y(2), ZN => L2_shift_L33_n_194);
  L2_shift_L33_g12997 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_177, A2 => L2_shift_L33_n_152, ZN => L2_shift_L33_n_319);
  L2_shift_L33_g12998 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_170, A2 => L2_shift_L33_n_149, ZN => L2_shift_L33_n_301);
  L2_shift_L33_g12999 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_177, A2 => L2_shift_L33_n_149, ZN => L2_shift_L33_n_305);
  L2_shift_L33_g13000 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_181, B1 => L2_shift_L33_n_149, ZN => L2_shift_L33_n_320);
  L2_shift_L33_g13001 : MAOI22D0BWP7T port map(A1 => L2_shift_L33_n_159, A2 => L2_shift_gg_pos_x(2), B1 => L2_shift_L33_n_159, B2 => L2_shift_gg_pos_x(2), ZN => L2_shift_L33_n_193);
  L2_shift_L33_g13002 : OA21D0BWP7T port map(A1 => L2_shift_L33_n_163, A2 => L2_shift_L33_n_147, B => L2_shift_L33_n_187, Z => L2_shift_L33_n_192);
  L2_shift_L33_g13003 : OA21D0BWP7T port map(A1 => L2_shift_L33_n_162, A2 => L2_shift_L33_n_146, B => L2_shift_L33_n_188, Z => L2_shift_L33_n_191);
  L2_shift_L33_g13004 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_178, B1 => L2_shift_L33_n_154, ZN => L2_shift_L33_n_310);
  L2_shift_L33_g13005 : AN3D1BWP7T port map(A1 => L2_shift_L33_n_153, A2 => L2_shift_L33_state(2), A3 => L2_shift_L33_state(0), Z => L2_shift_L33_n_299);
  L2_shift_L33_g13006 : AN3D1BWP7T port map(A1 => L2_shift_L33_n_153, A2 => L2_shift_L33_state(3), A3 => L2_shift_L33_state(0), Z => L2_shift_L33_n_309);
  L2_shift_L33_g13007 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_181, B1 => L2_shift_L33_n_154, ZN => L2_shift_L33_n_304);
  L2_shift_L33_g13008 : INVD1BWP7T port map(I => L2_shift_L33_n_182, ZN => L2_shift_L33_n_183);
  L2_shift_L33_g13009 : INVD1BWP7T port map(I => L2_shift_L33_n_179, ZN => L2_shift_L33_n_180);
  L2_shift_L33_g13010 : INVD0BWP7T port map(I => L2_shift_L33_n_177, ZN => L2_shift_L33_n_176);
  L2_shift_L33_g13011 : INR2XD0BWP7T port map(A1 => L2_shift_L33_n_159, B1 => L2_shift_L33_n_162, ZN => L2_shift_L33_n_190);
  L2_shift_L33_g13012 : OR2D1BWP7T port map(A1 => L2_shift_L33_n_159, A2 => L2_shift_L33_n_146, Z => L2_shift_L33_n_189);
  L2_shift_L33_g13013 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_162, A2 => L2_shift_L33_n_146, ZN => L2_shift_L33_n_188);
  L2_shift_L33_g13014 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_163, A2 => L2_shift_L33_n_147, ZN => L2_shift_L33_n_187);
  L2_shift_L33_g13015 : OR2D1BWP7T port map(A1 => L2_shift_L33_n_157, A2 => L2_shift_L33_n_147, Z => L2_shift_L33_n_186);
  L2_shift_L33_g13016 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_161, A2 => L2_shift_L33_n_154, ZN => L2_shift_L33_n_306);
  L2_shift_L33_g13017 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_161, B1 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_185);
  L2_shift_L33_g13018 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_155, A2 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_184);
  L2_shift_L33_g13019 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_294, B1 => L2_county(0), ZN => L2_shift_L33_n_293);
  L2_shift_L33_g13020 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_160, A2 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_182);
  L2_shift_L33_g13021 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_164, B1 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_181);
  L2_shift_L33_g13022 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_161, A2 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_179);
  L2_shift_L33_g13023 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_156, A2 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_178);
  L2_shift_L33_g13024 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_164, A2 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_177);
  L2_shift_L33_g13027 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(2), A2 => L2_shift_L33_n_146, B1 => xcoordinates_int(2), B2 => L2_shift_L33_n_146, ZN => L2_shift_L33_n_167);
  L2_shift_L33_g13028 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(2), A2 => L2_shift_L33_n_147, B1 => ycoordinates_int(2), B2 => L2_shift_L33_n_147, ZN => L2_shift_L33_n_166);
  L2_shift_L33_g13029 : CKXOR2D1BWP7T port map(A1 => xcoordinates_int(1), A2 => L2_shift_gg_pos_x(1), Z => L2_shift_L33_n_165);
  L2_shift_L33_g13030 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_144, A2 => L2_in_go_y_pos(1), B1 => L2_shift_L33_n_144, B2 => L2_in_go_y_pos(1), ZN => L2_shift_L33_n_175);
  L2_shift_L33_g13031 : AN2D0BWP7T port map(A1 => L2_shift_L33_n_294, A2 => L2_shift_L33_n_296, Z => L2_shift_L33_n_174);
  L2_shift_L33_g13032 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(0), A2 => L2_shift_gg_pos_y(0), Z => L2_shift_L33_n_173);
  L2_shift_L33_g13033 : CKXOR2D1BWP7T port map(A1 => xcoordinates_int(0), A2 => L2_shift_gg_pos_x(0), Z => L2_shift_L33_n_172);
  L2_shift_L33_g13034 : MAOI22D0BWP7T port map(A1 => ycoordinates_int(1), A2 => L2_shift_gg_pos_y(1), B1 => ycoordinates_int(1), B2 => L2_shift_gg_pos_y(1), ZN => L2_shift_L33_n_171);
  L2_shift_L33_g13035 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_53, A2 => L2_shift_L33_n_144, ZN => L2_shift_L33_n_297);
  L2_shift_L33_g13036 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_160, B1 => L2_shift_L33_state(0), ZN => L2_shift_L33_n_170);
  L2_shift_L33_g13037 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(4), A2 => L2_shift_gg_pos_x(4), B1 => xcoordinates_int(4), B2 => L2_shift_gg_pos_x(4), ZN => L2_shift_L33_n_169);
  L2_shift_L33_g13038 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(4), A2 => L2_shift_gg_pos_y(4), B1 => ycoordinates_int(4), B2 => L2_shift_gg_pos_y(4), ZN => L2_shift_L33_n_168);
  L2_shift_L33_g13039 : INVD0BWP7T port map(I => L2_shift_L33_n_53, ZN => L2_shift_L33_n_296);
  L2_shift_L33_g13040 : NR2D0BWP7T port map(A1 => L2_shift_L33_state(2), A2 => L2_shift_L33_state(3), ZN => L2_shift_L33_n_164);
  L2_shift_L33_g13041 : NR2XD0BWP7T port map(A1 => L2_shift_gg_pos_y(0), A2 => L2_shift_gg_pos_y(1), ZN => L2_shift_L33_n_163);
  L2_shift_L33_g13042 : NR2XD0BWP7T port map(A1 => L2_shift_gg_pos_x(0), A2 => L2_shift_gg_pos_x(1), ZN => L2_shift_L33_n_162);
  L2_shift_L33_g13043 : CKND2D1BWP7T port map(A1 => L2_shift_L33_state(2), A2 => L2_shift_L33_state(3), ZN => L2_shift_L33_n_161);
  L2_shift_L33_g13044 : IND2D1BWP7T port map(A1 => L2_shift_L33_state(3), B1 => L2_shift_L33_state(2), ZN => L2_shift_L33_n_160);
  L2_shift_L33_g13045 : ND2D1BWP7T port map(A1 => L2_shift_gg_pos_x(0), A2 => L2_shift_gg_pos_x(1), ZN => L2_shift_L33_n_159);
  L2_shift_L33_g13046 : NR2XD0BWP7T port map(A1 => L2_county(2), A2 => L2_in_go_y_pos(1), ZN => L2_shift_L33_n_53);
  L2_shift_L33_g13047 : INVD0BWP7T port map(I => L2_shift_L33_n_156, ZN => L2_shift_L33_n_155);
  L2_shift_L33_g13048 : INVD0BWP7T port map(I => L2_shift_L33_n_154, ZN => L2_shift_L33_n_153);
  L2_shift_L33_g13049 : INVD1BWP7T port map(I => L2_shift_L33_n_150, ZN => L2_shift_L33_n_149);
  L2_shift_L33_g13050 : ND2D1BWP7T port map(A1 => L2_shift_gg_pos_y(0), A2 => L2_shift_gg_pos_y(1), ZN => L2_shift_L33_n_157);
  L2_shift_L33_g13051 : IND2D1BWP7T port map(A1 => L2_shift_L33_state(2), B1 => L2_shift_L33_state(3), ZN => L2_shift_L33_n_156);
  L2_shift_L33_g13052 : CKND2D1BWP7T port map(A1 => L2_county(2), A2 => L2_in_go_y_pos(1), ZN => L2_shift_L33_n_294);
  L2_shift_L33_g13053 : CKND2D1BWP7T port map(A1 => L2_shift_L33_state(4), A2 => L2_shift_L33_state(1), ZN => L2_shift_L33_n_154);
  L2_shift_L33_g13054 : CKND2D1BWP7T port map(A1 => L2_shift_L33_n_145, A2 => L2_shift_L33_state(1), ZN => L2_shift_L33_n_152);
  L2_shift_L33_g13055 : IND2D1BWP7T port map(A1 => L2_shift_L33_state(1), B1 => L2_shift_L33_n_145, ZN => L2_shift_L33_n_151);
  L2_shift_L33_g13056 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_145, A2 => L2_shift_L33_state(1), ZN => L2_shift_L33_n_150);
  L2_shift_L33_g13060 : INVD0BWP7T port map(I => L2_county(2), ZN => L2_shift_L33_n_52);
  L2_shift_L33_g13062 : INVD1BWP7T port map(I => L2_shift_gg_pos_y(2), ZN => L2_shift_L33_n_147);
  L2_shift_L33_g13063 : INVD1BWP7T port map(I => L2_shift_gg_pos_x(2), ZN => L2_shift_L33_n_146);
  L2_shift_L33_g13065 : INVD1BWP7T port map(I => L2_county(0), ZN => L2_shift_L33_n_144);
  L2_shift_L33_g2 : CKXOR2D1BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_gg_pos_x(3), Z => L2_shift_L33_n_143);
  L2_shift_L33_g13066 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_gg_pos_y(3), Z => L2_shift_L33_n_142);
  L2_shift_L33_g10654 : AO211D0BWP7T port map(A1 => L2_pixel_array_to_shift(1), A2 => L2_shift_L33_n_65, B => L2_shift_L33_n_123, C => L2_shift_L33_n_139, Z => L2_shift_pixel_arr_out_shift_gg(0));
  L2_shift_L33_g10655 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_87, A2 => L2_shift_L33_n_55, B => L2_shift_L33_n_120, C => L2_shift_L33_n_136, ZN => L2_shift_pixel_arr_out_shift_gg(7));
  L2_shift_L33_g10656 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_75, A2 => L2_shift_L33_n_55, B => L2_shift_L33_n_119, C => L2_shift_L33_n_135, ZN => L2_shift_pixel_arr_out_shift_gg(6));
  L2_shift_L33_g10657 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_86, A2 => L2_shift_L33_n_55, B => L2_shift_L33_n_138, C => L2_shift_L33_n_116, ZN => L2_shift_pixel_arr_out_shift_gg(5));
  L2_shift_L33_g10658 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_85, A2 => L2_shift_L33_n_55, B => L2_shift_L33_n_141, C => L2_shift_L33_n_118, ZN => L2_shift_pixel_arr_out_shift_gg(3));
  L2_shift_L33_g10659 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_71, A2 => L2_shift_L33_n_55, B => L2_shift_L33_n_140, C => L2_shift_L33_n_117, ZN => L2_shift_pixel_arr_out_shift_gg(4));
  L2_shift_L33_g10660 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_67, A2 => L2_shift_L33_n_55, B => L2_shift_L33_n_137, C => L2_shift_L33_n_115, ZN => L2_shift_pixel_arr_out_shift_gg(2));
  L2_shift_L33_g10661 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_396, A2 => L2_shift_L33_n_55, B => L2_shift_L33_n_122, C => L2_shift_L33_n_114, ZN => L2_shift_pixel_arr_out_shift_gg(1));
  L2_shift_L33_g10662 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L33_n_68, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L33_n_65, C => L2_shift_L33_n_134, ZN => L2_shift_L33_n_141);
  L2_shift_L33_g10663 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(4), A2 => L2_shift_L33_n_131, B1 => L2_pixel_array_to_shift(5), B2 => L2_shift_L33_n_65, C => L2_shift_L33_n_106, ZN => L2_shift_L33_n_140);
  L2_shift_L33_g10664 : OAI22D0BWP7T port map(A1 => L2_shift_L33_n_49, A2 => L2_shift_L33_n_133, B1 => L2_shift_L33_n_51, B2 => L2_shift_L33_n_77, ZN => L2_shift_L33_n_139);
  L2_shift_L33_g10665 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L33_n_131, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L33_n_66, C => L2_shift_L33_n_103, ZN => L2_shift_L33_n_138);
  L2_shift_L33_g10666 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(2), A2 => L2_shift_L33_n_131, B1 => L2_pixel_array_to_shift(3), B2 => L2_shift_L33_n_65, C => L2_shift_L33_n_105, ZN => L2_shift_L33_n_137);
  L2_shift_L33_g10667 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L33_n_132, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L33_n_66, ZN => L2_shift_L33_n_136);
  L2_shift_L33_g10668 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(6), A2 => L2_shift_L33_n_131, B1 => L2_pixel_array_to_shift(7), B2 => L2_shift_L33_n_102, ZN => L2_shift_L33_n_135);
  L2_shift_L33_g10669 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L33_n_131, B1 => L2_shift_L33_n_66, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L33_n_134);
  L2_shift_L33_g10670 : AOI221D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_319, B1 => L2_shift_L33_n_394, B2 => L2_shift_L33_n_320, C => L2_shift_L33_n_131, ZN => L2_shift_L33_n_133);
  L2_shift_L33_g10671 : AO221D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_313, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_326, C => L2_shift_L33_n_131, Z => L2_shift_L33_n_132);
  L2_shift_L33_g10672 : INVD1BWP7T port map(I => L2_shift_L33_n_396, ZN => L2_shift_L33_n_131);
  L2_shift_L33_g10674 : IND4D0BWP7T port map(A1 => L2_shift_L33_n_283, B1 => L2_shift_L33_n_128, B2 => L2_shift_L33_n_127, B3 => L2_shift_L33_n_62, ZN => L2_shift_L33_n_129);
  L2_shift_L33_g10675 : AOI211XD0BWP7T port map(A1 => L2_shift_L33_n_289, A2 => L2_shift_L33_n_112, B => L2_shift_L33_n_126, C => L2_shift_L33_n_121, ZN => L2_shift_L33_n_128);
  L2_shift_L33_g10676 : AOI211XD0BWP7T port map(A1 => L2_shift_L33_n_290, A2 => L2_shift_L33_n_313, B => L2_shift_L33_n_124, C => L2_shift_L33_n_91, ZN => L2_shift_L33_n_127);
  L2_shift_L33_g10677 : IND4D0BWP7T port map(A1 => L2_shift_L33_n_288, B1 => L2_shift_L33_n_82, B2 => L2_shift_L33_n_83, B3 => L2_shift_L33_n_125, ZN => L2_shift_L33_n_126);
  L2_shift_L33_g10678 : AO211D0BWP7T port map(A1 => L2_shift_L33_n_113, A2 => L2_shift_L33_n_387, B => L2_shift_gg_pos_reset, C => L2_shift_L33_n_327, Z => L2_shift_shift_clock_reset_gg);
  L2_shift_L33_g10679 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_395, A2 => L2_shift_L33_n_111, B1 => L2_shift_L33_n_290, B2 => L2_shift_L33_n_92, ZN => L2_shift_L33_n_125);
  L2_shift_L33_g10680 : OAI222D0BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_99, B1 => L2_shift_L33_n_88, B2 => L2_shift_L33_n_393, C1 => L2_shift_L33_n_95, C2 => L2_shift_L33_n_61, ZN => L2_shift_L33_n_124);
  L2_shift_L33_g10681 : OAI221D0BWP7T port map(A1 => L2_shift_L33_n_57, A2 => L2_shift_L33_n_76, B1 => L2_shift_L33_n_74, B2 => L2_shift_L33_n_50, C => L2_shift_L33_n_104, ZN => L2_shift_L33_n_123);
  L2_shift_L33_g10682 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L33_n_68, B1 => L2_pixel_array_to_shift(2), B2 => L2_shift_L33_n_65, C => L2_shift_L33_n_110, ZN => L2_shift_L33_n_122);
  L2_shift_L33_g10683 : AOI21D0BWP7T port map(A1 => L2_shift_L33_n_89, A2 => L2_shift_L33_n_63, B => L2_shift_L33_n_298, ZN => L2_shift_L33_n_121);
  L2_shift_L33_g10684 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L33_n_84, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L33_n_70, C => L2_shift_L33_n_108, ZN => L2_shift_L33_n_120);
  L2_shift_L33_g10685 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L33_n_66, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L33_n_84, C => L2_shift_L33_n_107, ZN => L2_shift_L33_n_119);
  L2_shift_L33_g10686 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L33_n_98, B1 => L2_shift_L33_n_51, B2 => L2_shift_L33_n_73, ZN => L2_shift_L33_n_118);
  L2_shift_L33_g10687 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L33_n_96, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L33_n_68, ZN => L2_shift_L33_n_117);
  L2_shift_L33_g10688 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L33_n_97, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L33_n_65, ZN => L2_shift_L33_n_116);
  L2_shift_L33_g10689 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L33_n_101, B1 => L2_shift_L33_n_51, B2 => L2_shift_L33_n_74, ZN => L2_shift_L33_n_115);
  L2_shift_L33_g10690 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L33_n_100, B1 => L2_shift_L33_n_51, B2 => L2_shift_L33_n_76, ZN => L2_shift_L33_n_114);
  L2_shift_L33_g10691 : OR2D1BWP7T port map(A1 => L2_shift_L33_n_391, A2 => L2_shift_L33_n_94, Z => L2_shift_L33_n_113);
  L2_shift_L33_g10692 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => xcoordinates_int(0), Z => L2_shift_gg_pos_x_new(0));
  L2_shift_L33_g10693 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => xcoordinates_int(3), Z => L2_shift_gg_pos_x_new(3));
  L2_shift_L33_g10694 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => ycoordinates_int(4), Z => L2_shift_gg_pos_y_new(4));
  L2_shift_L33_g10695 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => ycoordinates_int(3), Z => L2_shift_gg_pos_y_new(3));
  L2_shift_L33_g10696 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_302, B1 => L2_shift_L33_n_93, ZN => L2_shift_L33_n_112);
  L2_shift_L33_g10697 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => ycoordinates_int(2), Z => L2_shift_gg_pos_y_new(2));
  L2_shift_L33_g10698 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => xcoordinates_int(4), Z => L2_shift_gg_pos_x_new(4));
  L2_shift_L33_g10699 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => ycoordinates_int(1), Z => L2_shift_gg_pos_y_new(1));
  L2_shift_L33_g10700 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_322, B1 => L2_shift_L33_n_90, ZN => L2_shift_L33_n_111);
  L2_shift_L33_g10701 : OAI22D0BWP7T port map(A1 => L2_shift_L33_n_57, A2 => L2_shift_L33_n_74, B1 => L2_shift_L33_n_50, B2 => L2_shift_L33_n_73, ZN => L2_shift_L33_n_110);
  L2_shift_L33_g10702 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => xcoordinates_int(1), Z => L2_shift_gg_pos_x_new(1));
  L2_shift_L33_g10703 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => xcoordinates_int(2), Z => L2_shift_gg_pos_x_new(2));
  L2_shift_L33_g10704 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_80, B => L2_shift_L33_n_81, ZN => L2_shift_L33_n_109);
  L2_shift_L33_g10705 : OAI22D0BWP7T port map(A1 => L2_shift_L33_n_58, A2 => L2_shift_L33_n_86, B1 => L2_shift_L33_n_56, B2 => L2_shift_L33_n_75, ZN => L2_shift_L33_n_108);
  L2_shift_L33_g10706 : AN2D0BWP7T port map(A1 => L2_shift_gg_pos_load, A2 => ycoordinates_int(0), Z => L2_shift_gg_pos_y_new(0));
  L2_shift_L33_g10707 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_56, A2 => L2_shift_L33_n_86, B1 => L2_pixel_array_to_shift(3), B2 => L2_shift_L33_n_70, ZN => L2_shift_L33_n_107);
  L2_shift_L33_g10708 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L33_n_66, B1 => L2_shift_L33_n_84, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L33_n_106);
  L2_shift_L33_g10709 : OAI22D0BWP7T port map(A1 => L2_shift_L33_n_57, A2 => L2_shift_L33_n_73, B1 => L2_shift_L33_n_50, B2 => L2_shift_L33_n_69, ZN => L2_shift_L33_n_105);
  L2_shift_L33_g10710 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L33_n_72, B1 => L2_pixel_array_to_shift(2), B2 => L2_shift_L33_n_68, ZN => L2_shift_L33_n_104);
  L2_shift_L33_g10711 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L33_n_84, B1 => L2_shift_L33_n_70, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L33_n_103);
  L2_shift_L33_g10712 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_87, A2 => L2_shift_L33_n_64, ZN => L2_shift_L33_n_102);
  L2_shift_L33_g10713 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_85, A2 => L2_shift_L33_n_76, ZN => L2_shift_L33_n_101);
  L2_shift_L33_g10714 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_67, A2 => L2_shift_L33_n_77, ZN => L2_shift_L33_n_100);
  L2_shift_L33_g10715 : AOI221D0BWP7T port map(A1 => L2_shift_L33_n_293, A2 => L2_shift_L33_n_306, B1 => L2_shift_L33_n_307, B2 => L2_shift_L33_n_294, C => L2_shift_L33_n_79, ZN => L2_shift_L33_n_99);
  L2_shift_L33_g10716 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_71, A2 => L2_shift_L33_n_74, ZN => L2_shift_L33_n_98);
  L2_shift_L33_g10717 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_75, A2 => L2_shift_L33_n_69, ZN => L2_shift_L33_n_97);
  L2_shift_L33_g10718 : ND2D1BWP7T port map(A1 => L2_shift_L33_n_86, A2 => L2_shift_L33_n_73, ZN => L2_shift_L33_n_96);
  L2_shift_L33_g10719 : INR2XD0BWP7T port map(A1 => L2_shift_L33_n_387, B1 => L2_shift_L33_n_391, ZN => L2_shift_gg_pos_load);
  L2_shift_L33_g10720 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_308, A2 => L2_shift_L33_n_307, A3 => L2_shift_L33_n_309, A4 => L2_shift_L33_n_306, ZN => L2_shift_L33_n_95);
  L2_shift_L33_g10721 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_393, A3 => L2_shift_L33_n_328, A4 => L2_shift_L33_n_394, ZN => L2_shift_L33_n_94);
  L2_shift_L33_g10722 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_301, A2 => L2_shift_L33_n_305, A3 => L2_shift_L33_n_304, A4 => L2_shift_L33_n_303, ZN => L2_shift_L33_n_93);
  L2_shift_L33_g10723 : OR4D1BWP7T port map(A1 => L2_shift_L33_n_316, A2 => L2_shift_L33_n_315, A3 => L2_shift_L33_n_317, A4 => L2_shift_L33_n_314, Z => L2_shift_L33_n_92);
  L2_shift_L33_g10724 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_61, A2 => L2_shift_L33_n_78, ZN => L2_shift_L33_n_91);
  L2_shift_L33_g10725 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_326, A2 => L2_shift_L33_n_325, A3 => L2_shift_L33_n_324, A4 => L2_shift_L33_n_323, ZN => L2_shift_L33_n_90);
  L2_shift_L33_g10726 : AOI222D0BWP7T port map(A1 => L2_shift_L33_n_301, A2 => L2_shift_L33_n_59, B1 => L2_shift_L33_n_305, B2 => L2_shift_L33_n_293, C1 => L2_shift_L33_n_302, C2 => L2_shift_L33_n_52, ZN => L2_shift_L33_n_89);
  L2_shift_L33_g10727 : AOI222D0BWP7T port map(A1 => L2_shift_L33_n_310, A2 => L2_shift_L33_n_59, B1 => L2_shift_L33_n_312, B2 => L2_shift_L33_n_54, C1 => L2_shift_L33_n_311, C2 => L2_shift_L33_n_53, ZN => L2_shift_L33_n_88);
  L2_shift_L33_g10728 : INVD1BWP7T port map(I => L2_shift_L33_n_85, ZN => L2_shift_L33_n_84);
  L2_shift_L33_g10729 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_319, A2 => L2_shift_L33_n_318, B => L2_shift_L33_n_290, ZN => L2_shift_L33_n_83);
  L2_shift_L33_g10730 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_320, A2 => L2_shift_L33_n_321, B => L2_shift_L33_n_395, ZN => L2_shift_L33_n_82);
  L2_shift_L33_g10731 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_300, A2 => L2_shift_L33_n_299, B => L2_shift_L33_n_289, ZN => L2_shift_L33_n_81);
  L2_shift_L33_g10732 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_299, A2 => L2_shift_L33_n_54, B1 => L2_shift_L33_n_300, B2 => L2_shift_L33_n_53, ZN => L2_shift_L33_n_80);
  L2_shift_L33_g10733 : AO22D0BWP7T port map(A1 => L2_shift_L33_n_309, A2 => L2_shift_L33_n_52, B1 => L2_shift_L33_n_279, B2 => L2_shift_L33_n_308, Z => L2_shift_L33_n_79);
  L2_shift_L33_g10734 : NR3D0BWP7T port map(A1 => L2_shift_L33_n_310, A2 => L2_shift_L33_n_312, A3 => L2_shift_L33_n_311, ZN => L2_shift_L33_n_78);
  L2_shift_L33_g10735 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_314, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_325, ZN => L2_shift_L33_n_87);
  L2_shift_L33_g10736 : IND3D1BWP7T port map(A1 => cell_type_int(2), B1 => cell_type_int(1), B2 => cell_type_int(0), ZN => L2_shift_L33_n_391);
  L2_shift_L33_g10737 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_316, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_323, ZN => L2_shift_L33_n_86);
  L2_shift_L33_g10738 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_318, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_321, ZN => L2_shift_L33_n_85);
  L2_shift_L33_g10739 : INVD0BWP7T port map(I => L2_shift_L33_n_73, ZN => L2_shift_L33_n_72);
  L2_shift_L33_g10740 : INVD1BWP7T port map(I => L2_shift_L33_n_71, ZN => L2_shift_L33_n_70);
  L2_shift_L33_g10741 : INVD1BWP7T port map(I => L2_shift_L33_n_69, ZN => L2_shift_L33_n_68);
  L2_shift_L33_g10742 : INVD1BWP7T port map(I => L2_shift_L33_n_67, ZN => L2_shift_L33_n_66);
  L2_shift_L33_g10743 : INVD1BWP7T port map(I => L2_shift_L33_n_64, ZN => L2_shift_L33_n_65);
  L2_shift_L33_g10744 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_303, A2 => L2_shift_L33_n_279, B1 => L2_shift_L33_n_304, B2 => L2_shift_L33_n_294, ZN => L2_shift_L33_n_63);
  L2_shift_L33_g10745 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_280, A2 => L2_shift_L33_n_286, A3 => L2_shift_L33_n_281, A4 => L2_shift_L33_n_282, ZN => L2_shift_L33_n_62);
  L2_shift_L33_g10746 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_318, B1 => L2_shift_L33_n_394, B2 => L2_shift_L33_n_321, ZN => L2_shift_L33_n_77);
  L2_shift_L33_g10747 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_317, B1 => L2_shift_L33_n_394, B2 => L2_shift_L33_n_322, ZN => L2_shift_L33_n_76);
  L2_shift_L33_g10748 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_315, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_324, ZN => L2_shift_L33_n_75);
  L2_shift_L33_g10749 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_316, B1 => L2_shift_L33_n_394, B2 => L2_shift_L33_n_323, ZN => L2_shift_L33_n_74);
  L2_shift_L33_g10750 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_315, B1 => L2_shift_L33_n_394, B2 => L2_shift_L33_n_324, ZN => L2_shift_L33_n_73);
  L2_shift_L33_g10751 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_317, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_322, ZN => L2_shift_L33_n_71);
  L2_shift_L33_g10752 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_314, B1 => L2_shift_L33_n_394, B2 => L2_shift_L33_n_325, ZN => L2_shift_L33_n_69);
  L2_shift_L33_g10753 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_319, B1 => L2_shift_L33_n_298, B2 => L2_shift_L33_n_320, ZN => L2_shift_L33_n_67);
  L2_shift_L33_g10754 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_298, A2 => L2_shift_L33_n_313, B1 => L2_shift_L33_n_394, B2 => L2_shift_L33_n_326, ZN => L2_shift_L33_n_64);
  L2_shift_L33_g10755 : OR2D1BWP7T port map(A1 => L2_shift_L33_n_393, A2 => L2_shift_L33_n_298, Z => L2_shift_L33_n_61);
  L2_shift_L33_g10757 : INVD0BWP7T port map(I => L2_shift_L33_n_295, ZN => L2_shift_L33_n_59);
  L2_shift_L33_g10758 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(3), ZN => L2_shift_L33_n_58);
  L2_shift_L33_g10759 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(5), ZN => L2_shift_L33_n_57);
  L2_shift_L33_g10760 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(2), ZN => L2_shift_L33_n_56);
  L2_shift_L33_g10761 : INVD1BWP7T port map(I => L2_pixel_array_to_shift(1), ZN => L2_shift_L33_n_55);
  L2_shift_L33_g10762 : INVD0BWP7T port map(I => L2_shift_L33_n_297, ZN => L2_shift_L33_n_54);
  L2_shift_L33_g10765 : INVD1BWP7T port map(I => L2_pixel_array_to_shift(6), ZN => L2_shift_L33_n_51);
  L2_shift_L33_g10766 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(4), ZN => L2_shift_L33_n_50);
  L2_shift_L33_g10767 : CKND1BWP7T port map(I => L2_pixel_array_to_shift(7), ZN => L2_shift_L33_n_49);
  L2_shift_L33_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L33_n_48, Q => L2_shift_L33_state(0));
  L2_shift_L33_g10068 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_47, A2 => L2_shift_L33_n_6, A3 => L2_shift_L33_n_15, A4 => L2_shift_L33_n_0, ZN => L2_shift_L33_n_48);
  L2_shift_L33_state_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L33_n_46, Q => L2_shift_L33_state(3));
  L2_shift_L33_g10070 : OAI211D1BWP7T port map(A1 => L2_shift_L33_n_2, A2 => L2_shift_L33_n_5, B => L2_shift_L33_n_18, C => L2_shift_L33_n_45, ZN => L2_shift_L33_n_47);
  L2_shift_L33_g10071 : ND4D0BWP7T port map(A1 => L2_shift_L33_n_26, A2 => L2_shift_L33_n_25, A3 => L2_shift_L33_n_41, A4 => L2_shift_L33_n_27, ZN => L2_shift_L33_n_46);
  L2_shift_L33_g10072 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_42, A2 => L2_shift_shift_pulse_gg, B1 => L2_shift_L33_n_32, B2 => L2_shift_shift_pulse_gg, ZN => L2_shift_L33_n_45);
  L2_shift_L33_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L33_n_44, Q => L2_shift_L33_state(1));
  L2_shift_L33_g10075 : IND4D0BWP7T port map(A1 => L2_shift_L33_n_15, B1 => L2_shift_L33_n_12, B2 => L2_shift_L33_n_26, B3 => L2_shift_L33_n_39, ZN => L2_shift_L33_n_44);
  L2_shift_L33_g10076 : IND4D0BWP7T port map(A1 => L2_shift_L33_n_38, B1 => L2_shift_L33_n_16, B2 => L2_shift_L33_n_17, B3 => L2_shift_L33_n_12, ZN => L2_shift_L33_n_43);
  L2_shift_L33_g10077 : IINR4D0BWP7T port map(A1 => L2_shift_L33_n_37, A2 => L2_shift_L33_n_5, B1 => L2_shift_L33_n_313, B2 => L2_shift_L33_n_387, ZN => L2_shift_L33_n_42);
  L2_shift_L33_state_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L33_n_40, Q => L2_shift_L33_state(2));
  L2_shift_L33_g10079 : AOI221D0BWP7T port map(A1 => L2_shift_L33_n_36, A2 => L2_shift_L33_n_1, B1 => L2_shift_L33_n_313, B2 => L2_shift_L33_n_4, C => L2_shift_L33_n_20, ZN => L2_shift_L33_n_41);
  L2_shift_L33_g10080 : IND4D0BWP7T port map(A1 => L2_shift_L33_n_29, B1 => L2_shift_L33_n_27, B2 => L2_shift_L33_n_31, B3 => L2_shift_L33_n_33, ZN => L2_shift_L33_n_40);
  L2_shift_L33_g10081 : NR3D0BWP7T port map(A1 => L2_shift_L33_n_24, A2 => L2_shift_L33_n_34, A3 => L2_shift_L33_n_29, ZN => L2_shift_L33_n_39);
  L2_shift_L33_g10082 : ND4D0BWP7T port map(A1 => L2_shift_L33_n_30, A2 => L2_shift_L33_n_25, A3 => L2_shift_L33_n_31, A4 => L2_shift_L33_n_19, ZN => L2_shift_L33_n_38);
  L2_shift_L33_g10083 : INR4D0BWP7T port map(A1 => L2_shift_L33_n_32, B1 => L2_shift_L33_n_299, B2 => L2_shift_L33_n_327, B3 => L2_shift_gg_pos_reset, ZN => L2_shift_L33_n_37);
  L2_shift_L33_g10084 : IND2D1BWP7T port map(A1 => L2_shift_L33_n_325, B1 => L2_shift_L33_n_35, ZN => L2_shift_L33_n_36);
  L2_shift_L33_g10085 : NR4D0BWP7T port map(A1 => L2_shift_L33_n_22, A2 => L2_shift_L33_n_310, A3 => L2_shift_L33_n_311, A4 => L2_shift_L33_n_307, ZN => L2_shift_L33_n_35);
  L2_shift_L33_g10086 : AO221D0BWP7T port map(A1 => L2_shift_L33_n_28, A2 => L2_shift_shift_pulse_gg, B1 => L2_shift_L33_n_23, B2 => L2_shift_L33_n_2, C => L2_shift_L33_n_21, Z => L2_shift_L33_n_34);
  L2_shift_L33_g10087 : AOI222D0BWP7T port map(A1 => L2_shift_L33_n_23, A2 => L2_shift_shift_pulse_gg, B1 => L2_shift_L33_n_8, B2 => L2_shift_L33_n_1, C1 => L2_shift_L33_n_315, C2 => L2_shift_L33_n_4, ZN => L2_shift_L33_n_33);
  L2_shift_L33_g10088 : NR2XD0BWP7T port map(A1 => L2_shift_L33_n_28, A2 => L2_shift_L33_n_23, ZN => L2_shift_L33_n_32);
  L2_shift_L33_g10089 : AOI222D0BWP7T port map(A1 => L2_shift_L33_n_11, A2 => L2_shift_L33_n_393, B1 => L2_shift_L33_n_320, B2 => L2_shift_L33_n_4, C1 => L2_shift_L33_n_9, C2 => L2_shift_L33_n_1, ZN => L2_shift_L33_n_30);
  L2_shift_L33_g10090 : AOI211XD0BWP7T port map(A1 => L2_shift_L33_n_302, A2 => L2_shift_L33_n_1, B => L2_shift_L33_n_13, C => L2_shift_L33_n_20, ZN => L2_shift_L33_n_31);
  L2_shift_L33_g10091 : IOA21D1BWP7T port map(A1 => L2_shift_L33_n_316, A2 => L2_shift_L33_n_1, B => L2_shift_L33_n_19, ZN => L2_shift_L33_n_29);
  L2_shift_L33_g10092 : IND3D1BWP7T port map(A1 => L2_shift_L33_n_13, B1 => L2_shift_L33_n_10, B2 => L2_shift_L33_n_17, ZN => L2_shift_L33_n_28);
  L2_shift_L33_g10093 : MAOI22D0BWP7T port map(A1 => L2_shift_L33_n_321, A2 => L2_shift_L33_n_4, B1 => L2_shift_L33_n_14, B2 => L2_shift_L33_n_0, ZN => L2_shift_L33_n_27);
  L2_shift_L33_g10094 : MOAI22D0BWP7T port map(A1 => L2_shift_L33_n_5, A2 => L2_shift_L33_n_3, B1 => L2_shift_L33_n_11, B2 => L2_shift_L33_n_394, ZN => L2_shift_L33_n_24);
  L2_shift_L33_g10095 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_11, A2 => L2_shift_L33_n_287, B1 => L2_shift_L33_n_326, B2 => L2_shift_L33_n_1, ZN => L2_shift_L33_n_26);
  L2_shift_L33_g10096 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_11, A2 => L2_shift_L33_n_328, B1 => L2_shift_L33_n_312, B2 => L2_shift_L33_n_1, ZN => L2_shift_L33_n_25);
  L2_shift_L33_g10097 : AO211D0BWP7T port map(A1 => L2_shift_L33_n_315, A2 => L2_shift_shift_pulse_gg, B => L2_shift_L33_n_314, C => L2_shift_L33_n_309, Z => L2_shift_L33_n_22);
  L2_shift_L33_g10098 : OA21D0BWP7T port map(A1 => L2_shift_L33_n_6, A2 => L2_shift_L33_n_322, B => L2_shift_L33_n_1, Z => L2_shift_L33_n_21);
  L2_shift_L33_g10099 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_7, A2 => L2_shift_L33_n_0, B => L2_shift_L33_n_16, ZN => L2_shift_L33_n_23);
  L2_shift_L33_g10100 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_287, A2 => L2_shift_L33_n_328, B => L2_shift_L33_n_11, ZN => L2_shift_L33_n_18);
  L2_shift_L33_g10101 : AO21D0BWP7T port map(A1 => L2_shift_L33_n_308, A2 => L2_shift_L33_n_1, B => L2_shift_L33_n_15, Z => L2_shift_L33_n_20);
  L2_shift_L33_g10102 : AOI22D0BWP7T port map(A1 => L2_shift_L33_n_299, A2 => L2_shift_L33_n_4, B1 => L2_shift_L33_n_300, B2 => L2_shift_L33_n_1, ZN => L2_shift_L33_n_19);
  L2_shift_L33_g10103 : NR3D0BWP7T port map(A1 => L2_shift_L33_n_322, A2 => L2_shift_L33_n_323, A3 => L2_shift_L33_n_324, ZN => L2_shift_L33_n_14);
  L2_shift_L33_g10104 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_311, A2 => L2_shift_L33_n_305, B => L2_shift_L33_n_1, ZN => L2_shift_L33_n_17);
  L2_shift_L33_g10105 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_309, A2 => L2_shift_L33_n_303, B => L2_shift_L33_n_1, ZN => L2_shift_L33_n_16);
  L2_shift_L33_g10106 : AN2D1BWP7T port map(A1 => L2_shift_L33_n_306, A2 => L2_shift_L33_n_4, Z => L2_shift_L33_n_15);
  L2_shift_L33_g10107 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_317, A2 => L2_shift_L33_n_323, B => L2_shift_L33_n_1, ZN => L2_shift_L33_n_10);
  L2_shift_L33_g10108 : OA21D0BWP7T port map(A1 => L2_shift_L33_n_301, A2 => L2_shift_L33_n_307, B => L2_shift_L33_n_1, Z => L2_shift_L33_n_13);
  L2_shift_L33_g10109 : OAI21D0BWP7T port map(A1 => L2_shift_L33_n_310, A2 => L2_shift_L33_n_304, B => L2_shift_L33_n_1, ZN => L2_shift_L33_n_12);
  L2_shift_L33_g10110 : INR3D0BWP7T port map(A1 => L2_shift_L33_n_387, B1 => L2_shift_L33_n_0, B2 => L2_shift_L33_n_391, ZN => L2_shift_L33_n_11);
  L2_shift_L33_g10111 : AN2D0BWP7T port map(A1 => L2_shift_L33_n_321, A2 => L2_shift_shift_pulse_gg, Z => L2_shift_L33_n_9);
  L2_shift_L33_g10112 : OR2D1BWP7T port map(A1 => L2_shift_L33_n_317, A2 => L2_shift_L33_n_318, Z => L2_shift_L33_n_8);
  L2_shift_L33_g10113 : NR2D0BWP7T port map(A1 => L2_shift_L33_n_325, A2 => L2_shift_L33_n_319, ZN => L2_shift_L33_n_7);
  L2_shift_L33_g10114 : INVD0BWP7T port map(I => L2_shift_L33_n_4, ZN => L2_shift_L33_n_3);
  L2_shift_L33_g10115 : INR2D1BWP7T port map(A1 => L2_shift_L33_n_327, B1 => L2_calc_start_internal, ZN => L2_shift_L33_n_6);
  L2_shift_L33_g10116 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_315, A2 => L2_shift_L33_n_321, ZN => L2_shift_L33_n_5);
  L2_shift_L33_g10117 : NR2D1BWP7T port map(A1 => L2_shift_L33_n_0, A2 => L2_shift_shift_pulse_gg, ZN => L2_shift_L33_n_4);
  L2_shift_L33_g10118 : INVD0BWP7T port map(I => L2_shift_shift_pulse_gg, ZN => L2_shift_L33_n_2);
  L2_shift_L33_drc_bufs10120 : INVD1BWP7T port map(I => L2_shift_L33_n_1, ZN => L2_shift_L33_n_0);
  L2_shift_L33_drc_bufs10121 : INVD0BWP7T port map(I => reset, ZN => L2_shift_L33_n_1);
  L2_shift_L33_g13067 : NR2D0BWP7T port map(A1 => L2_shift_L33_n_394, A2 => L2_shift_L33_n_298, ZN => L2_shift_L33_n_395);
  L2_shift_L33_state_reg_4 : DFD1BWP7T port map(CP => clk, D => L2_shift_L33_n_43, Q => L2_shift_L33_state(4), QN => L2_shift_L33_n_145);
  L2_shift_L33_g13070 : INR4D0BWP7T port map(A1 => L2_shift_L33_n_257, B1 => L2_shift_L33_n_129, B2 => L2_shift_L33_n_285, B3 => L2_shift_L33_n_109, ZN => L2_shift_L33_n_396);
  L2_shift_L21_shift_sync_gr_reg : DFQD0BWP7T port map(CP => clk, D => L2_shift_L21_n_9, Q => L2_shift_shift_pulse_gr);
  L2_shift_L21_g174 : INR4D0BWP7T port map(A1 => L2_calc_start_internal, B1 => L2_shift_L21_count_internal(0), B2 => L2_shift_L21_n_8, B3 => L2_shift_shift_clock_reset_gr, ZN => L2_shift_L21_n_9);
  L2_shift_L21_g175 : IND2D1BWP7T port map(A1 => L2_shift_L21_count_internal(1), B1 => L2_shift_L21_count_internal(2), ZN => L2_shift_L21_n_8);
  L2_shift_L21_count_internal_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L21_n_7, Q => L2_shift_L21_count_internal(2));
  L2_shift_L21_count_internal_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L21_n_6, Q => L2_shift_L21_count_internal(1));
  L2_shift_L21_g244 : AO22D0BWP7T port map(A1 => L2_shift_L21_n_3, A2 => L2_shift_L21_n_4, B1 => L2_shift_L21_count_internal(2), B2 => L2_shift_L21_n_1, Z => L2_shift_L21_n_7);
  L2_shift_L21_g246 : AO22D0BWP7T port map(A1 => L2_shift_L21_n_3, A2 => L2_shift_L21_n_2, B1 => L2_shift_L21_count_internal(1), B2 => L2_shift_L21_n_1, Z => L2_shift_L21_n_6);
  L2_shift_L21_g247 : AO22D0BWP7T port map(A1 => L2_shift_L21_n_3, A2 => L2_shift_L21_n_10, B1 => L2_shift_L21_count_internal(0), B2 => L2_shift_L21_n_1, Z => L2_shift_L21_n_5);
  L2_shift_L21_g248 : MOAI22D0BWP7T port map(A1 => L2_shift_L21_n_0, A2 => L2_shift_L21_count_internal(2), B1 => L2_shift_L21_n_0, B2 => L2_shift_L21_count_internal(2), ZN => L2_shift_L21_n_4);
  L2_shift_L21_g249 : NR3D0BWP7T port map(A1 => L2_shift_L21_n_9, A2 => L2_shift_L21_n_1, A3 => L2_shift_shift_clock_reset_gr, ZN => L2_shift_L21_n_3);
  L2_shift_L21_g250 : MOAI22D0BWP7T port map(A1 => L2_shift_L21_n_10, A2 => L2_shift_L21_count_internal(1), B1 => L2_shift_L21_n_10, B2 => L2_shift_L21_count_internal(1), ZN => L2_shift_L21_n_2);
  L2_shift_L21_g251 : NR2XD0BWP7T port map(A1 => L2_shift_shift_clock_reset_gr, A2 => L2_calc_start_internal, ZN => L2_shift_L21_n_1);
  L2_shift_L21_g252 : ND2D1BWP7T port map(A1 => L2_shift_L21_count_internal(1), A2 => L2_shift_L21_count_internal(0), ZN => L2_shift_L21_n_0);
  L2_shift_L21_count_internal_reg_0 : DFD1BWP7T port map(CP => clk, D => L2_shift_L21_n_5, Q => L2_shift_L21_count_internal(0), QN => L2_shift_L21_n_10);
  L2_shift_L23_g17610 : IND4D0BWP7T port map(A1 => L2_shift_L23_n_260, B1 => L2_shift_L23_n_399, B2 => L2_shift_L23_n_269, B3 => L2_shift_L23_n_279, ZN => L2_shift_y_pos_out_shift_gr(2));
  L2_shift_L23_g17611 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_275, A2 => L2_county(0), B => L2_shift_L23_n_281, ZN => L2_shift_y_pos_out_shift_gr(0));
  L2_shift_L23_g17612 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_183, A2 => L2_shift_L23_n_272, B => L2_shift_L23_n_280, C => L2_shift_L23_n_271, ZN => L2_shift_y_pos_out_shift_gr(1));
  L2_shift_L23_g17613 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_278, A2 => L2_shift_L23_n_268, B => L2_county(0), ZN => L2_shift_L23_n_281);
  L2_shift_L23_g17614 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_278, A2 => L2_in_go_y_pos(1), B1 => L2_shift_L23_n_263, B2 => L2_shift_L23_n_183, ZN => L2_shift_L23_n_280);
  L2_shift_L23_g17615 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_277, A2 => L2_county(2), B1 => L2_shift_L23_n_331, B2 => L2_shift_L23_n_305, ZN => L2_shift_L23_n_279);
  L2_shift_L23_g17616 : OR2D1BWP7T port map(A1 => L2_shift_L23_n_277, A2 => L2_shift_L23_n_286, Z => L2_shift_L23_n_278);
  L2_shift_L23_g17617 : IINR4D0BWP7T port map(A1 => L2_shift_L23_n_276, A2 => L2_shift_L23_n_259, B1 => L2_shift_L23_n_285, B2 => L2_shift_L23_n_286, ZN => L2_shift_L23_n_277);
  L2_shift_L23_g17618 : AN2D0BWP7T port map(A1 => cell_type_int(2), A2 => L2_shift_L23_n_274, Z => L2_shift_cell_state_out_shift_gr(2));
  L2_shift_L23_g17619 : AN2D0BWP7T port map(A1 => cell_type_int(0), A2 => L2_shift_L23_n_274, Z => L2_shift_cell_state_out_shift_gr(0));
  L2_shift_L23_g17620 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_268, A2 => L2_shift_L23_n_263, A3 => L2_shift_L23_n_289, A4 => L2_shift_L23_n_283, ZN => L2_shift_L23_n_276);
  L2_shift_L23_g17621 : IOA21D1BWP7T port map(A1 => L2_shift_L23_n_267, A2 => L2_shift_L23_n_301, B => L2_shift_L23_n_273, ZN => L2_shift_cell_state_out_shift_gr(1));
  L2_shift_L23_g17622 : INR2XD0BWP7T port map(A1 => L2_shift_L23_n_272, B1 => L2_shift_L23_n_263, ZN => L2_shift_L23_n_275);
  L2_shift_L23_g17623 : IAO21D0BWP7T port map(A1 => L2_shift_L23_n_265, A2 => L2_shift_L23_n_267, B => cell_type_int(1), ZN => L2_shift_L23_n_273);
  L2_shift_L23_g17624 : IOA21D1BWP7T port map(A1 => L2_shift_L23_n_267, A2 => L2_shift_L23_n_228, B => L2_shift_L23_n_264, ZN => L2_shift_L23_n_274);
  L2_shift_L23_g17625 : AO21D0BWP7T port map(A1 => L2_shift_L23_n_262, A2 => L2_shift_L23_n_256, B => L2_in_go_y_pos(1), Z => L2_shift_L23_n_271);
  L2_shift_L23_g17626 : INR3D0BWP7T port map(A1 => L2_shift_L23_n_259, B1 => L2_shift_L23_n_285, B2 => L2_shift_L23_n_261, ZN => L2_shift_L23_n_272);
  L2_shift_L23_g17628 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_257, A2 => L2_shift_L23_n_209, B1 => L2_shift_L23_n_261, B2 => L2_shift_L23_n_208, ZN => L2_shift_L23_n_269);
  L2_shift_L23_g17629 : IND3D0BWP7T port map(A1 => L2_shift_L23_n_284, B1 => L2_shift_L23_n_256, B2 => L2_shift_L23_n_255, ZN => L2_shift_L23_n_268);
  L2_shift_L23_g17631 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_397, A2 => L2_shift_L23_n_221, B1 => L2_shift_L23_n_396, B2 => L2_shift_L23_n_196, ZN => L2_shift_L23_n_267);
  L2_shift_L23_g17632 : INVD1BWP7T port map(I => L2_shift_L23_n_264, ZN => L2_shift_L23_n_265);
  L2_shift_L23_g17633 : AOI221D0BWP7T port map(A1 => L2_shift_L23_n_292, A2 => L2_shift_L23_n_226, B1 => L2_shift_L23_n_293, B2 => L2_shift_L23_n_220, C => L2_shift_L23_n_291, ZN => L2_shift_L23_n_264);
  L2_shift_L23_g17634 : IND2D1BWP7T port map(A1 => L2_shift_L23_n_257, B1 => L2_shift_L23_n_254, ZN => L2_shift_L23_n_263);
  L2_shift_L23_g17635 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_254, A2 => L2_shift_L23_n_209, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_312, ZN => L2_shift_L23_n_260);
  L2_shift_L23_g17636 : AOI21D0BWP7T port map(A1 => L2_shift_L23_n_247, A2 => L2_shift_L23_n_59, B => L2_shift_L23_n_288, ZN => L2_shift_L23_n_262);
  L2_shift_L23_g17637 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_244, A2 => L2_shift_L23_n_300, B => L2_shift_L23_n_258, ZN => L2_shift_L23_n_261);
  L2_shift_L23_g17638 : INVD0BWP7T port map(I => L2_shift_L23_n_289, ZN => L2_shift_L23_n_258);
  L2_shift_L23_g17639 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_246, A2 => L2_shift_L23_n_282, ZN => L2_shift_L23_n_259);
  L2_shift_L23_g17640 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_248, A2 => L2_shift_L23_n_282, ZN => L2_shift_L23_n_285);
  L2_shift_L23_g17641 : INR2XD0BWP7T port map(A1 => L2_shift_L23_n_300, B1 => L2_shift_L23_n_251, ZN => L2_shift_L23_n_289);
  L2_shift_L23_g17642 : INVD0BWP7T port map(I => L2_shift_L23_n_288, ZN => L2_shift_L23_n_255);
  L2_shift_L23_g17643 : AOI211XD0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L23_n_219, B => L2_shift_L23_n_252, C => L2_shift_L23_n_230, ZN => L2_shift_L23_n_397);
  L2_shift_L23_g17644 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_240, A2 => L2_shift_L23_n_298, B => L2_shift_L23_n_253, ZN => L2_shift_L23_n_257);
  L2_shift_L23_g17645 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_250, A2 => L2_shift_L23_n_297, ZN => L2_shift_L23_n_256);
  L2_shift_L23_g17646 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_249, A2 => L2_shift_L23_n_59, ZN => L2_shift_L23_n_288);
  L2_shift_L23_g17648 : ND4D0BWP7T port map(A1 => L2_shift_L23_n_218, A2 => L2_shift_L23_n_236, A3 => L2_shift_L23_n_203, A4 => L2_shift_L23_n_177, ZN => L2_shift_L23_n_252);
  L2_shift_L23_g17649 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_241, A2 => L2_shift_L23_n_296, ZN => L2_shift_L23_n_254);
  L2_shift_L23_g17650 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_245, A2 => L2_shift_L23_n_298, ZN => L2_shift_L23_n_253);
  L2_shift_L23_g17651 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_243, A2 => L2_shift_L23_n_297, ZN => L2_shift_L23_n_284);
  L2_shift_L23_g17652 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_239, A2 => L2_shift_L23_n_296, ZN => L2_shift_L23_n_283);
  L2_shift_L23_g17653 : CKAN2D1BWP7T port map(A1 => L2_shift_L23_n_242, A2 => L2_county(2), Z => L2_shift_L23_n_286);
  L2_shift_L23_g17654 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_237, A2 => L2_shift_L23_n_186, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_302, ZN => L2_shift_L23_n_251);
  L2_shift_L23_g17655 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_238, A2 => L2_shift_L23_n_170, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_310, ZN => L2_shift_L23_n_250);
  L2_shift_L23_g17656 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_237, A2 => L2_shift_L23_n_188, B1 => L2_shift_L23_n_234, B2 => L2_shift_L23_n_185, ZN => L2_shift_L23_n_249);
  L2_shift_L23_g17657 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_237, A2 => L2_shift_L23_n_187, B1 => L2_shift_L23_n_234, B2 => L2_shift_L23_n_168, ZN => L2_shift_L23_n_248);
  L2_shift_L23_g17658 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_238, A2 => L2_shift_L23_n_184, B1 => L2_shift_L23_n_233, B2 => L2_shift_L23_n_189, ZN => L2_shift_L23_n_247);
  L2_shift_L23_g17659 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_238, A2 => L2_shift_L23_n_169, B1 => L2_shift_L23_n_233, B2 => L2_shift_L23_n_143, ZN => L2_shift_L23_n_246);
  L2_shift_L23_g17660 : AO22D0BWP7T port map(A1 => L2_shift_L23_n_396, A2 => L2_shift_L23_n_313, B1 => L2_shift_L23_n_304, B2 => L2_shift_L23_n_301, Z => L2_shift_L23_n_245);
  L2_shift_L23_g17661 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_331, A2 => L2_shift_L23_n_302, B1 => L2_shift_L23_n_232, B2 => L2_shift_L23_n_186, ZN => L2_shift_L23_n_244);
  L2_shift_L23_g17662 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_396, A2 => L2_shift_L23_n_310, B1 => L2_shift_L23_n_234, B2 => L2_shift_L23_n_171, ZN => L2_shift_L23_n_243);
  L2_shift_L23_g17663 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_301, ZN => L2_shift_L23_n_293);
  L2_shift_L23_g17664 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_233, A2 => L2_shift_L23_n_184, B1 => L2_shift_L23_n_396, B2 => L2_shift_L23_n_312, ZN => L2_shift_L23_n_242);
  L2_shift_L23_g17665 : AO22D0BWP7T port map(A1 => L2_shift_L23_n_331, A2 => L2_shift_L23_n_308, B1 => L2_shift_L23_n_309, B2 => L2_shift_L23_n_301, Z => L2_shift_L23_n_241);
  L2_shift_L23_g17666 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_331, A2 => L2_shift_L23_n_304, B1 => L2_shift_L23_n_234, B2 => L2_shift_L23_n_186, ZN => L2_shift_L23_n_240);
  L2_shift_L23_g17667 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_396, A2 => L2_shift_L23_n_309, B1 => L2_shift_L23_n_232, B2 => L2_shift_L23_n_168, ZN => L2_shift_L23_n_239);
  L2_shift_L23_g17668 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_331, A2 => L2_shift_L23_n_301, ZN => L2_shift_L23_n_292);
  L2_shift_L23_g17669 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_331, A2 => L2_shift_L23_n_151, ZN => L2_shift_L23_n_238);
  L2_shift_L23_g17670 : AOI211XD0BWP7T port map(A1 => xcoordinates_int(2), A2 => L2_shift_L23_n_197, B => L2_shift_L23_n_235, C => L2_shift_L23_n_214, ZN => L2_shift_L23_n_290);
  L2_shift_L23_g17671 : CKAN2D1BWP7T port map(A1 => L2_shift_L23_n_396, A2 => L2_shift_L23_n_161, Z => L2_shift_L23_n_237);
  L2_shift_L23_g17672 : AOI221D0BWP7T port map(A1 => L2_shift_L23_n_173, A2 => L2_shift_L23_n_210, B1 => xcoordinates_int(2), B2 => L2_shift_L23_n_198, C => L2_shift_L23_n_231, ZN => L2_shift_L23_n_236);
  L2_shift_L23_g17673 : NR3D0BWP7T port map(A1 => L2_shift_L23_n_227, A2 => L2_shift_L23_n_225, A3 => L2_shift_L23_n_204, ZN => L2_shift_L23_n_331);
  L2_shift_L23_g17674 : IND4D0BWP7T port map(A1 => L2_shift_L23_n_203, B1 => L2_shift_L23_n_177, B2 => L2_shift_L23_n_224, B3 => L2_shift_L23_n_218, ZN => L2_shift_L23_n_235);
  L2_shift_L23_g17675 : NR3D0BWP7T port map(A1 => L2_shift_L23_n_229, A2 => L2_shift_L23_n_225, A3 => L2_shift_L23_n_216, ZN => L2_shift_L23_n_396);
  L2_shift_L23_g17676 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_228, A2 => L2_shift_L23_n_152, ZN => L2_shift_L23_n_234);
  L2_shift_L23_g17677 : CKND1BWP7T port map(I => L2_shift_L23_n_233, ZN => L2_shift_L23_n_232);
  L2_shift_L23_g17678 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_173, A2 => L2_shift_L23_n_210, B1 => xcoordinates_int(2), B2 => L2_shift_L23_n_198, ZN => L2_shift_L23_n_231);
  L2_shift_L23_g17679 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_161, ZN => L2_shift_L23_n_233);
  L2_shift_L23_g17680 : NR2D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L23_n_219, ZN => L2_shift_L23_n_230);
  L2_shift_L23_g17681 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_194, A2 => L2_shift_L23_n_207, B => L2_shift_L23_n_223, C => L2_shift_L23_n_204, ZN => L2_shift_L23_n_229);
  L2_shift_L23_g17682 : INVD0BWP7T port map(I => L2_shift_L23_n_301, ZN => L2_shift_L23_n_228);
  L2_shift_L23_g17683 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_222, A2 => L2_shift_L23_n_215, B1 => L2_shift_L23_n_212, B2 => L2_shift_L23_n_158, ZN => L2_shift_L23_n_227);
  L2_shift_L23_g17684 : AN3D1BWP7T port map(A1 => L2_shift_L23_n_218, A2 => L2_shift_L23_n_211, A3 => L2_shift_L23_n_173, Z => L2_shift_L23_n_301);
  L2_shift_L23_g17685 : OR4D1BWP7T port map(A1 => L2_shift_L23_n_302, A2 => L2_shift_L23_n_307, A3 => L2_shift_L23_n_304, A4 => L2_shift_L23_n_205, Z => L2_shift_L23_n_226);
  L2_shift_L23_g17686 : AOI211XD0BWP7T port map(A1 => L2_shift_L23_n_180, A2 => L2_shift_L23_n_195, B => L2_shift_L23_n_217, C => L2_shift_L23_n_201, ZN => L2_shift_L23_n_224);
  L2_shift_L23_g17687 : ND3D0BWP7T port map(A1 => L2_shift_L23_n_211, A2 => L2_shift_L23_n_178, A3 => L2_shift_L23_n_173, ZN => L2_shift_L23_n_225);
  L2_shift_L23_g17688 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_200, A2 => L2_shift_L23_n_166, B => L2_shift_L23_n_194, ZN => L2_shift_L23_n_223);
  L2_shift_L23_g17689 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_142, A2 => L2_shift_L23_n_166, B => L2_shift_gr_pos_y(2), ZN => L2_shift_L23_n_222);
  L2_shift_L23_g17690 : AOI211XD0BWP7T port map(A1 => L2_shift_L23_n_191, A2 => L2_shift_L23_n_160, B => L2_shift_L23_n_202, C => L2_shift_L23_n_323, ZN => L2_shift_L23_n_221);
  L2_shift_L23_g17691 : AO211D0BWP7T port map(A1 => L2_shift_L23_n_164, A2 => L2_shift_L23_n_162, B => L2_shift_L23_n_206, C => L2_shift_L23_n_322, Z => L2_shift_L23_n_220);
  L2_shift_L23_g17692 : AOI211D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L23_n_149, B => L2_shift_L23_n_172, C => L2_shift_L23_n_195, ZN => L2_shift_L23_n_217);
  L2_shift_L23_g17693 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(2), A2 => L2_shift_L23_n_199, B1 => ycoordinates_int(2), B2 => L2_shift_L23_n_199, ZN => L2_shift_L23_n_216);
  L2_shift_L23_g17694 : NR3D0BWP7T port map(A1 => L2_shift_L23_n_213, A2 => L2_shift_L23_n_179, A3 => L2_shift_L23_n_158, ZN => L2_shift_L23_n_215);
  L2_shift_L23_g17695 : AOI21D0BWP7T port map(A1 => L2_shift_L23_n_192, A2 => L2_shift_gr_pos_x(3), B => L2_shift_L23_n_210, ZN => L2_shift_L23_n_219);
  L2_shift_L23_g17696 : INR3D0BWP7T port map(A1 => L2_shift_L23_n_212, B1 => L2_shift_L23_n_178, B2 => L2_shift_L23_n_175, ZN => L2_shift_L23_n_218);
  L2_shift_L23_g17697 : NR2D0BWP7T port map(A1 => xcoordinates_int(2), A2 => L2_shift_L23_n_197, ZN => L2_shift_L23_n_214);
  L2_shift_L23_g17698 : NR2D0BWP7T port map(A1 => L2_shift_L23_n_207, A2 => L2_shift_gr_pos_y(2), ZN => L2_shift_L23_n_213);
  L2_shift_L23_g17699 : CKAN2D1BWP7T port map(A1 => L2_shift_L23_n_207, A2 => L2_shift_L23_n_179, Z => L2_shift_L23_n_212);
  L2_shift_L23_g17700 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_180, A2 => L2_shift_L23_n_177, A3 => L2_shift_L23_n_176, A4 => L2_shift_L23_n_167, ZN => L2_shift_L23_n_211);
  L2_shift_L23_g17701 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_192, A2 => L2_shift_gr_pos_x(3), ZN => L2_shift_L23_n_210);
  L2_shift_L23_g17702 : IAO21D0BWP7T port map(A1 => L2_shift_L23_n_185, A2 => L2_shift_L23_n_190, B => L2_shift_L23_state(4), ZN => L2_shift_L23_n_206);
  L2_shift_L23_g17703 : OA21D0BWP7T port map(A1 => L2_shift_L23_n_185, A2 => L2_shift_L23_n_168, B => L2_shift_L23_state(4), Z => L2_shift_L23_n_205);
  L2_shift_L23_g17704 : OAI211D1BWP7T port map(A1 => L2_county(0), A2 => L2_county(2), B => L2_shift_L23_n_296, C => L2_shift_L23_n_299, ZN => L2_shift_L23_n_209);
  L2_shift_L23_g17705 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_144, A2 => L2_shift_L23_n_58, B => L2_shift_L23_n_300, C => L2_shift_L23_n_297, ZN => L2_shift_L23_n_208);
  L2_shift_L23_g17706 : AO21D0BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(0), B => L2_county(2), Z => L2_shift_L23_n_298);
  L2_shift_L23_g17707 : OAI21D0BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(0), B => L2_county(2), ZN => L2_shift_L23_n_282);
  L2_shift_L23_g17708 : AOI211XD0BWP7T port map(A1 => L2_shift_L23_n_150, A2 => L2_shift_gr_pos_y(3), B => L2_shift_L23_n_174, C => L2_shift_L23_n_159, ZN => L2_shift_L23_n_207);
  L2_shift_L23_g17709 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_143, A2 => L2_shift_L23_state(4), B1 => L2_shift_L23_n_164, B2 => L2_shift_L23_n_163, ZN => L2_shift_L23_n_202);
  L2_shift_L23_g17710 : IAO21D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L23_n_149, B => L2_shift_L23_n_173, ZN => L2_shift_L23_n_201);
  L2_shift_L23_g17712 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_174, A2 => L2_shift_L23_n_150, B1 => L2_shift_L23_n_174, B2 => L2_shift_gr_pos_y(3), ZN => L2_shift_L23_n_200);
  L2_shift_L23_g17713 : CKXOR2D1BWP7T port map(A1 => L2_shift_L23_n_175, A2 => L2_shift_gr_pos_y(0), Z => L2_shift_L23_n_204);
  L2_shift_L23_g17714 : AO21D0BWP7T port map(A1 => L2_shift_L23_n_171, A2 => L2_shift_L23_n_145, B => L2_shift_L23_n_390, Z => L2_shift_L23_n_291);
  L2_shift_L23_g17715 : MAOI22D0BWP7T port map(A1 => L2_shift_L23_n_176, A2 => L2_shift_gr_pos_x(0), B1 => L2_shift_L23_n_176, B2 => L2_shift_gr_pos_x(0), ZN => L2_shift_L23_n_203);
  L2_shift_L23_g17716 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_162, B1 => L2_shift_L23_n_170, ZN => L2_shift_gr_pos_reset);
  L2_shift_L23_g17717 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_190, A2 => L2_shift_L23_n_162, Z => L2_shift_L23_n_320);
  L2_shift_L23_g17718 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_190, A2 => L2_shift_L23_n_163, Z => L2_shift_L23_n_318);
  L2_shift_L23_g17719 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_191, A2 => L2_shift_L23_state(1), Z => L2_shift_L23_n_324);
  L2_shift_L23_g17720 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_189, A2 => L2_shift_L23_n_160, ZN => L2_shift_L23_n_314);
  L2_shift_L23_g17721 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_163, B1 => L2_shift_L23_n_170, ZN => L2_shift_L23_n_330);
  L2_shift_L23_g17722 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_163, B1 => L2_shift_L23_n_189, ZN => L2_shift_L23_n_328);
  L2_shift_L23_g17723 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_162, B1 => L2_shift_L23_n_189, ZN => L2_shift_L23_n_316);
  L2_shift_L23_g17724 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_186, A2 => L2_shift_L23_n_162, Z => L2_shift_L23_n_317);
  L2_shift_L23_g17725 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_162, B1 => L2_shift_L23_n_184, ZN => L2_shift_L23_n_321);
  L2_shift_L23_g17726 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_162, B1 => L2_shift_L23_n_169, ZN => L2_shift_L23_n_390);
  L2_shift_L23_g17727 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_170, A2 => L2_shift_L23_n_160, ZN => L2_shift_L23_n_323);
  L2_shift_L23_g17728 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_170, A2 => L2_shift_L23_n_152, ZN => L2_shift_L23_n_307);
  L2_shift_L23_g17729 : INR2XD0BWP7T port map(A1 => L2_shift_L23_state(2), B1 => L2_shift_L23_n_193, ZN => L2_shift_L23_n_309);
  L2_shift_L23_g17730 : INR2XD0BWP7T port map(A1 => L2_shift_L23_state(0), B1 => L2_shift_L23_n_193, ZN => L2_shift_L23_n_312);
  L2_shift_L23_g17731 : CKAN2D1BWP7T port map(A1 => L2_shift_L23_n_191, A2 => L2_shift_L23_state(4), Z => L2_shift_L23_n_310);
  L2_shift_L23_g17732 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_190, A2 => L2_shift_L23_n_161, Z => L2_shift_L23_n_304);
  L2_shift_L23_g17733 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_162, B1 => L2_shift_L23_n_143, ZN => L2_shift_L23_n_327);
  L2_shift_L23_g17734 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_143, A2 => L2_shift_L23_n_160, ZN => L2_shift_L23_n_311);
  L2_shift_L23_g17735 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_163, B1 => L2_shift_L23_n_143, ZN => L2_shift_L23_n_325);
  L2_shift_L23_g17736 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_186, B1 => L2_shift_L23_n_160, ZN => L2_shift_L23_n_315);
  L2_shift_L23_g17737 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_186, A2 => L2_shift_L23_n_163, Z => L2_shift_L23_n_329);
  L2_shift_L23_g17738 : OA21D0BWP7T port map(A1 => L2_shift_L23_n_160, A2 => L2_shift_L23_n_146, B => L2_shift_L23_n_193, Z => L2_shift_L23_n_196);
  L2_shift_L23_g17739 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_169, A2 => L2_shift_L23_n_152, ZN => L2_shift_L23_n_306);
  L2_shift_L23_g17740 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_184, A2 => L2_shift_L23_n_152, ZN => L2_shift_L23_n_303);
  L2_shift_L23_g17741 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_191, A2 => L2_shift_L23_n_162, Z => L2_shift_L23_n_326);
  L2_shift_L23_g17742 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_163, B1 => L2_shift_L23_n_184, ZN => L2_shift_L23_n_319);
  L2_shift_L23_g17743 : CKAN2D1BWP7T port map(A1 => L2_shift_L23_n_186, A2 => L2_shift_L23_n_151, Z => L2_shift_L23_n_313);
  L2_shift_L23_g17744 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_163, B1 => L2_shift_L23_n_169, ZN => L2_shift_L23_n_322);
  L2_shift_L23_g17745 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_184, A2 => L2_shift_L23_n_160, ZN => L2_shift_L23_n_305);
  L2_shift_L23_g17746 : AOI21D0BWP7T port map(A1 => L2_shift_L23_n_156, A2 => L2_shift_gr_pos_y(2), B => L2_shift_L23_n_194, ZN => L2_shift_L23_n_199);
  L2_shift_L23_g17747 : OA21D0BWP7T port map(A1 => L2_shift_L23_n_155, A2 => L2_shift_L23_n_148, B => L2_shift_L23_n_192, Z => L2_shift_L23_n_198);
  L2_shift_L23_g17748 : MAOI22D0BWP7T port map(A1 => L2_shift_L23_n_154, A2 => L2_shift_gr_pos_x(2), B1 => L2_shift_L23_n_154, B2 => L2_shift_gr_pos_x(2), ZN => L2_shift_L23_n_197);
  L2_shift_L23_g17749 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_169, A2 => L2_shift_L23_n_160, ZN => L2_shift_L23_n_308);
  L2_shift_L23_g17750 : CKND1BWP7T port map(I => L2_shift_L23_n_189, ZN => L2_shift_L23_n_188);
  L2_shift_L23_g17751 : INVD0BWP7T port map(I => L2_shift_L23_n_143, ZN => L2_shift_L23_n_187);
  L2_shift_L23_g17752 : INVD1BWP7T port map(I => L2_shift_L23_n_185, ZN => L2_shift_L23_n_184);
  L2_shift_L23_g17753 : OR2D1BWP7T port map(A1 => L2_shift_L23_n_154, A2 => L2_shift_L23_n_148, Z => L2_shift_L23_n_195);
  L2_shift_L23_g17754 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_156, A2 => L2_shift_gr_pos_y(2), ZN => L2_shift_L23_n_194);
  L2_shift_L23_g17755 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_151, A2 => L2_shift_L23_state(3), ZN => L2_shift_L23_n_193);
  L2_shift_L23_g17756 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_155, A2 => L2_shift_L23_n_148, ZN => L2_shift_L23_n_192);
  L2_shift_L23_g17757 : OR2D1BWP7T port map(A1 => L2_shift_L23_n_297, A2 => L2_shift_L23_n_144, Z => L2_shift_L23_n_296);
  L2_shift_L23_g17758 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_59, A2 => L2_shift_L23_n_144, ZN => L2_shift_L23_n_300);
  L2_shift_L23_g17759 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_165, A2 => L2_shift_L23_n_146, ZN => L2_shift_L23_n_191);
  L2_shift_L23_g17760 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_165, A2 => L2_shift_L23_n_152, ZN => L2_shift_L23_n_302);
  L2_shift_L23_g17761 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_165, A2 => L2_shift_L23_state(3), ZN => L2_shift_L23_n_190);
  L2_shift_L23_g17762 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_164, A2 => L2_shift_L23_state(0), ZN => L2_shift_L23_n_189);
  L2_shift_L23_g17764 : INR2XD0BWP7T port map(A1 => L2_shift_L23_n_164, B1 => L2_shift_L23_state(0), ZN => L2_shift_L23_n_186);
  L2_shift_L23_g17765 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_157, A2 => L2_shift_L23_state(3), ZN => L2_shift_L23_n_185);
  L2_shift_L23_g17766 : CKND1BWP7T port map(I => L2_shift_L23_n_181, ZN => L2_shift_L23_n_182);
  L2_shift_L23_g17767 : CKND1BWP7T port map(I => L2_shift_L23_n_173, ZN => L2_shift_L23_n_172);
  L2_shift_L23_g17768 : INVD1BWP7T port map(I => L2_shift_L23_n_171, ZN => L2_shift_L23_n_170);
  L2_shift_L23_g17769 : INVD0BWP7T port map(I => L2_shift_L23_n_169, ZN => L2_shift_L23_n_168);
  L2_shift_L23_g17770 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(2), A2 => L2_shift_L23_n_148, B1 => xcoordinates_int(2), B2 => L2_shift_L23_n_148, ZN => L2_shift_L23_n_167);
  L2_shift_L23_g17771 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_144, A2 => L2_in_go_y_pos(1), B1 => L2_shift_L23_n_144, B2 => L2_in_go_y_pos(1), ZN => L2_shift_L23_n_183);
  L2_shift_L23_g17772 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_299, A2 => L2_shift_L23_n_297, ZN => L2_shift_L23_n_181);
  L2_shift_L23_g17773 : MAOI22D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_gr_pos_x(3), B1 => xcoordinates_int(3), B2 => L2_shift_gr_pos_x(3), ZN => L2_shift_L23_n_180);
  L2_shift_L23_g17774 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(2), A2 => L2_shift_gr_pos_y(2), B1 => ycoordinates_int(2), B2 => L2_shift_gr_pos_y(2), ZN => L2_shift_L23_n_179);
  L2_shift_L23_g17775 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(0), A2 => L2_shift_gr_pos_y(0), Z => L2_shift_L23_n_178);
  L2_shift_L23_g17776 : CKXOR2D1BWP7T port map(A1 => xcoordinates_int(0), A2 => L2_shift_gr_pos_x(0), Z => L2_shift_L23_n_177);
  L2_shift_L23_g17777 : MAOI22D0BWP7T port map(A1 => xcoordinates_int(1), A2 => L2_shift_gr_pos_x(1), B1 => xcoordinates_int(1), B2 => L2_shift_gr_pos_x(1), ZN => L2_shift_L23_n_176);
  L2_shift_L23_g17778 : MAOI22D0BWP7T port map(A1 => ycoordinates_int(1), A2 => L2_shift_gr_pos_y(1), B1 => ycoordinates_int(1), B2 => L2_shift_gr_pos_y(1), ZN => L2_shift_L23_n_175);
  L2_shift_L23_g17779 : MAOI22D0BWP7T port map(A1 => ycoordinates_int(4), A2 => L2_shift_gr_pos_y(4), B1 => ycoordinates_int(4), B2 => L2_shift_gr_pos_y(4), ZN => L2_shift_L23_n_174);
  L2_shift_L23_g17780 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(4), A2 => L2_shift_gr_pos_x(4), B1 => xcoordinates_int(4), B2 => L2_shift_gr_pos_x(4), ZN => L2_shift_L23_n_173);
  L2_shift_L23_g17781 : NR3D0BWP7T port map(A1 => L2_shift_L23_state(3), A2 => L2_shift_L23_state(0), A3 => L2_shift_L23_state(2), ZN => L2_shift_L23_n_171);
  L2_shift_L23_g17782 : IND3D1BWP7T port map(A1 => L2_shift_L23_state(2), B1 => L2_shift_L23_state(0), B2 => L2_shift_L23_n_146, ZN => L2_shift_L23_n_169);
  L2_shift_L23_g17783 : INVD1BWP7T port map(I => L2_shift_L23_n_161, ZN => L2_shift_L23_n_160);
  L2_shift_L23_g17784 : NR2D0BWP7T port map(A1 => L2_shift_L23_n_150, A2 => L2_shift_gr_pos_y(3), ZN => L2_shift_L23_n_159);
  L2_shift_L23_g17785 : NR2D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_gr_pos_y(3), ZN => L2_shift_L23_n_166);
  L2_shift_L23_g17786 : CKND2D1BWP7T port map(A1 => L2_shift_L23_state(0), A2 => L2_shift_L23_state(2), ZN => L2_shift_L23_n_165);
  L2_shift_L23_g17787 : NR2XD0BWP7T port map(A1 => L2_shift_L23_n_146, A2 => L2_shift_L23_state(2), ZN => L2_shift_L23_n_164);
  L2_shift_L23_g17788 : INR2D1BWP7T port map(A1 => L2_shift_L23_state(1), B1 => L2_shift_L23_state(4), ZN => L2_shift_L23_n_163);
  L2_shift_L23_g17789 : NR2D1BWP7T port map(A1 => L2_shift_L23_state(4), A2 => L2_shift_L23_state(1), ZN => L2_shift_L23_n_162);
  L2_shift_L23_g17790 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_145, A2 => L2_shift_L23_state(1), ZN => L2_shift_L23_n_161);
  L2_shift_L23_g17792 : INVD1BWP7T port map(I => L2_shift_L23_n_59, ZN => L2_shift_L23_n_299);
  L2_shift_L23_g17793 : INVD1BWP7T port map(I => L2_shift_L23_n_152, ZN => L2_shift_L23_n_151);
  L2_shift_L23_g17794 : ND2D1BWP7T port map(A1 => L2_shift_gr_pos_y(0), A2 => L2_shift_gr_pos_y(1), ZN => L2_shift_L23_n_158);
  L2_shift_L23_g17795 : IND2D1BWP7T port map(A1 => L2_shift_L23_state(0), B1 => L2_shift_L23_state(2), ZN => L2_shift_L23_n_157);
  L2_shift_L23_g17796 : OR2D1BWP7T port map(A1 => L2_shift_gr_pos_y(0), A2 => L2_shift_gr_pos_y(1), Z => L2_shift_L23_n_156);
  L2_shift_L23_g17797 : NR2XD0BWP7T port map(A1 => L2_shift_gr_pos_x(1), A2 => L2_shift_gr_pos_x(0), ZN => L2_shift_L23_n_155);
  L2_shift_L23_g17798 : ND2D1BWP7T port map(A1 => L2_shift_gr_pos_x(1), A2 => L2_shift_gr_pos_x(0), ZN => L2_shift_L23_n_154);
  L2_shift_L23_g17799 : NR2D1BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(2), ZN => L2_shift_L23_n_59);
  L2_shift_L23_g17800 : CKND2D1BWP7T port map(A1 => L2_county(2), A2 => L2_in_go_y_pos(1), ZN => L2_shift_L23_n_297);
  L2_shift_L23_g17801 : CKND2D1BWP7T port map(A1 => L2_shift_L23_state(4), A2 => L2_shift_L23_state(1), ZN => L2_shift_L23_n_152);
  L2_shift_L23_g17802 : INVD0BWP7T port map(I => ycoordinates_int(3), ZN => L2_shift_L23_n_150);
  L2_shift_L23_g17803 : INVD0BWP7T port map(I => L2_shift_gr_pos_x(3), ZN => L2_shift_L23_n_149);
  L2_shift_L23_g17804 : INVD1BWP7T port map(I => L2_shift_gr_pos_x(2), ZN => L2_shift_L23_n_148);
  L2_shift_L23_g17809 : INVD1BWP7T port map(I => L2_county(0), ZN => L2_shift_L23_n_144);
  L2_shift_L23_g2 : IND2D1BWP7T port map(A1 => L2_shift_L23_n_157, B1 => L2_shift_L23_state(3), ZN => L2_shift_L23_n_143);
  L2_shift_L23_g17810 : MUX2D0BWP7T port map(I0 => L2_shift_gr_pos_y(3), I1 => ycoordinates_int(3), S => L2_shift_L23_n_174, Z => L2_shift_L23_n_142);
  L2_shift_L23_g10634 : AO211D0BWP7T port map(A1 => L2_pixel_array_to_shift(1), A2 => L2_shift_L23_n_68, B => L2_shift_L23_n_120, C => L2_shift_L23_n_139, Z => L2_shift_pixel_arr_out_shift_gr(0));
  L2_shift_L23_g10635 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_77, A2 => L2_shift_L23_n_56, B => L2_shift_L23_n_119, C => L2_shift_L23_n_136, ZN => L2_shift_pixel_arr_out_shift_gr(7));
  L2_shift_L23_g10636 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_76, A2 => L2_shift_L23_n_56, B => L2_shift_L23_n_118, C => L2_shift_L23_n_135, ZN => L2_shift_pixel_arr_out_shift_gr(6));
  L2_shift_L23_g10637 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_75, A2 => L2_shift_L23_n_56, B => L2_shift_L23_n_138, C => L2_shift_L23_n_117, ZN => L2_shift_pixel_arr_out_shift_gr(5));
  L2_shift_L23_g10638 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_86, A2 => L2_shift_L23_n_56, B => L2_shift_L23_n_141, C => L2_shift_L23_n_115, ZN => L2_shift_pixel_arr_out_shift_gr(3));
  L2_shift_L23_g10639 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_72, A2 => L2_shift_L23_n_56, B => L2_shift_L23_n_140, C => L2_shift_L23_n_116, ZN => L2_shift_pixel_arr_out_shift_gr(4));
  L2_shift_L23_g10640 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_66, A2 => L2_shift_L23_n_56, B => L2_shift_L23_n_137, C => L2_shift_L23_n_114, ZN => L2_shift_pixel_arr_out_shift_gr(2));
  L2_shift_L23_g10641 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_398, A2 => L2_shift_L23_n_56, B => L2_shift_L23_n_123, C => L2_shift_L23_n_113, ZN => L2_shift_pixel_arr_out_shift_gr(1));
  L2_shift_L23_g10642 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L23_n_69, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L23_n_68, C => L2_shift_L23_n_134, ZN => L2_shift_L23_n_141);
  L2_shift_L23_g10643 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(4), A2 => L2_shift_L23_n_131, B1 => L2_pixel_array_to_shift(5), B2 => L2_shift_L23_n_68, C => L2_shift_L23_n_106, ZN => L2_shift_L23_n_140);
  L2_shift_L23_g10644 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_51, A2 => L2_shift_L23_n_133, B1 => L2_shift_L23_n_57, B2 => L2_shift_L23_n_78, ZN => L2_shift_L23_n_139);
  L2_shift_L23_g10645 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L23_n_131, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L23_n_65, C => L2_shift_L23_n_103, ZN => L2_shift_L23_n_138);
  L2_shift_L23_g10646 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(2), A2 => L2_shift_L23_n_131, B1 => L2_pixel_array_to_shift(3), B2 => L2_shift_L23_n_68, C => L2_shift_L23_n_105, ZN => L2_shift_L23_n_137);
  L2_shift_L23_g10647 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L23_n_132, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L23_n_65, ZN => L2_shift_L23_n_136);
  L2_shift_L23_g10648 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(6), A2 => L2_shift_L23_n_131, B1 => L2_pixel_array_to_shift(7), B2 => L2_shift_L23_n_98, ZN => L2_shift_L23_n_135);
  L2_shift_L23_g10649 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L23_n_131, B1 => L2_shift_L23_n_65, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L23_n_134);
  L2_shift_L23_g10650 : AOI221D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_322, B1 => L2_shift_L23_n_397, B2 => L2_shift_L23_n_323, C => L2_shift_L23_n_131, ZN => L2_shift_L23_n_133);
  L2_shift_L23_g10651 : AO221D0BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_316, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_329, C => L2_shift_L23_n_131, Z => L2_shift_L23_n_132);
  L2_shift_L23_g10652 : INVD1BWP7T port map(I => L2_shift_L23_n_398, ZN => L2_shift_L23_n_131);
  L2_shift_L23_g10654 : IND4D0BWP7T port map(A1 => L2_shift_L23_n_286, B1 => L2_shift_L23_n_128, B2 => L2_shift_L23_n_126, B3 => L2_shift_L23_n_63, ZN => L2_shift_L23_n_129);
  L2_shift_L23_g10655 : AOI211XD0BWP7T port map(A1 => L2_shift_L23_n_292, A2 => L2_shift_L23_n_111, B => L2_shift_L23_n_127, C => L2_shift_L23_n_121, ZN => L2_shift_L23_n_128);
  L2_shift_L23_g10656 : IND4D0BWP7T port map(A1 => L2_shift_L23_n_291, B1 => L2_shift_L23_n_82, B2 => L2_shift_L23_n_122, B3 => L2_shift_L23_n_125, ZN => L2_shift_L23_n_127);
  L2_shift_L23_g10657 : AOI211XD0BWP7T port map(A1 => L2_shift_L23_n_293, A2 => L2_shift_L23_n_316, B => L2_shift_L23_n_124, C => L2_shift_L23_n_95, ZN => L2_shift_L23_n_126);
  L2_shift_L23_g10658 : OAI31D0BWP7T port map(A1 => L2_shift_L23_n_321, A2 => L2_shift_L23_n_322, A3 => L2_shift_L23_n_91, B => L2_shift_L23_n_293, ZN => L2_shift_L23_n_125);
  L2_shift_L23_g10659 : AO211D0BWP7T port map(A1 => L2_shift_L23_n_112, A2 => L2_shift_L23_n_390, B => L2_shift_gr_pos_reset, C => L2_shift_L23_n_330, Z => L2_shift_shift_clock_reset_gr);
  L2_shift_L23_g10660 : OAI222D0BWP7T port map(A1 => L2_shift_L23_n_396, A2 => L2_shift_L23_n_92, B1 => L2_shift_L23_n_89, B2 => L2_shift_L23_n_396, C1 => L2_shift_L23_n_96, C2 => L2_shift_L23_n_62, ZN => L2_shift_L23_n_124);
  L2_shift_L23_g10661 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L23_n_69, B1 => L2_pixel_array_to_shift(2), B2 => L2_shift_L23_n_68, C => L2_shift_L23_n_108, ZN => L2_shift_L23_n_123);
  L2_shift_L23_g10662 : OAI31D0BWP7T port map(A1 => L2_shift_L23_n_326, A2 => L2_shift_L23_n_325, A3 => L2_shift_L23_n_83, B => L2_shift_L23_n_61, ZN => L2_shift_L23_n_122);
  L2_shift_L23_g10663 : AOI21D0BWP7T port map(A1 => L2_shift_L23_n_90, A2 => L2_shift_L23_n_64, B => L2_shift_L23_n_301, ZN => L2_shift_L23_n_121);
  L2_shift_L23_g10664 : OAI221D0BWP7T port map(A1 => L2_shift_L23_n_49, A2 => L2_shift_L23_n_88, B1 => L2_shift_L23_n_87, B2 => L2_shift_L23_n_50, C => L2_shift_L23_n_104, ZN => L2_shift_L23_n_120);
  L2_shift_L23_g10665 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L23_n_85, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L23_n_71, C => L2_shift_L23_n_109, ZN => L2_shift_L23_n_119);
  L2_shift_L23_g10666 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L23_n_65, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L23_n_85, C => L2_shift_L23_n_107, ZN => L2_shift_L23_n_118);
  L2_shift_L23_g10667 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L23_n_97, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L23_n_68, ZN => L2_shift_L23_n_117);
  L2_shift_L23_g10668 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L23_n_102, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L23_n_69, ZN => L2_shift_L23_n_116);
  L2_shift_L23_g10669 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L23_n_99, B1 => L2_shift_L23_n_57, B2 => L2_shift_L23_n_74, ZN => L2_shift_L23_n_115);
  L2_shift_L23_g10670 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L23_n_101, B1 => L2_shift_L23_n_57, B2 => L2_shift_L23_n_87, ZN => L2_shift_L23_n_114);
  L2_shift_L23_g10671 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L23_n_100, B1 => L2_shift_L23_n_57, B2 => L2_shift_L23_n_88, ZN => L2_shift_L23_n_113);
  L2_shift_L23_g10672 : OR2D1BWP7T port map(A1 => L2_shift_L23_n_394, A2 => L2_shift_L23_n_94, Z => L2_shift_L23_n_112);
  L2_shift_L23_g10673 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => xcoordinates_int(0), Z => L2_shift_gr_pos_x_new(0));
  L2_shift_L23_g10674 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => xcoordinates_int(3), Z => L2_shift_gr_pos_x_new(3));
  L2_shift_L23_g10675 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => ycoordinates_int(4), Z => L2_shift_gr_pos_y_new(4));
  L2_shift_L23_g10676 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => ycoordinates_int(3), Z => L2_shift_gr_pos_y_new(3));
  L2_shift_L23_g10677 : IND2D1BWP7T port map(A1 => L2_shift_L23_n_305, B1 => L2_shift_L23_n_93, ZN => L2_shift_L23_n_111);
  L2_shift_L23_g10678 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => ycoordinates_int(2), Z => L2_shift_gr_pos_y_new(2));
  L2_shift_L23_g10679 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => ycoordinates_int(1), Z => L2_shift_gr_pos_y_new(1));
  L2_shift_L23_g10680 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => xcoordinates_int(4), Z => L2_shift_gr_pos_x_new(4));
  L2_shift_L23_g10681 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => ycoordinates_int(0), Z => L2_shift_gr_pos_y_new(0));
  L2_shift_L23_g10682 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => xcoordinates_int(2), Z => L2_shift_gr_pos_x_new(2));
  L2_shift_L23_g10683 : AN2D0BWP7T port map(A1 => L2_shift_gr_pos_load, A2 => xcoordinates_int(1), Z => L2_shift_gr_pos_x_new(1));
  L2_shift_L23_g10684 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_80, B => L2_shift_L23_n_81, ZN => L2_shift_L23_n_110);
  L2_shift_L23_g10685 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_54, A2 => L2_shift_L23_n_75, B1 => L2_shift_L23_n_55, B2 => L2_shift_L23_n_76, ZN => L2_shift_L23_n_109);
  L2_shift_L23_g10686 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_49, A2 => L2_shift_L23_n_87, B1 => L2_shift_L23_n_50, B2 => L2_shift_L23_n_74, ZN => L2_shift_L23_n_108);
  L2_shift_L23_g10687 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_55, A2 => L2_shift_L23_n_75, B1 => L2_pixel_array_to_shift(3), B2 => L2_shift_L23_n_71, ZN => L2_shift_L23_n_107);
  L2_shift_L23_g10688 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L23_n_65, B1 => L2_shift_L23_n_85, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L23_n_106);
  L2_shift_L23_g10689 : OAI22D0BWP7T port map(A1 => L2_shift_L23_n_49, A2 => L2_shift_L23_n_74, B1 => L2_shift_L23_n_50, B2 => L2_shift_L23_n_70, ZN => L2_shift_L23_n_105);
  L2_shift_L23_g10690 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L23_n_73, B1 => L2_pixel_array_to_shift(2), B2 => L2_shift_L23_n_69, ZN => L2_shift_L23_n_104);
  L2_shift_L23_g10691 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L23_n_85, B1 => L2_shift_L23_n_71, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L23_n_103);
  L2_shift_L23_g10692 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_75, A2 => L2_shift_L23_n_74, ZN => L2_shift_L23_n_102);
  L2_shift_L23_g10693 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_86, A2 => L2_shift_L23_n_88, ZN => L2_shift_L23_n_101);
  L2_shift_L23_g10694 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_66, A2 => L2_shift_L23_n_78, ZN => L2_shift_L23_n_100);
  L2_shift_L23_g10695 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_72, A2 => L2_shift_L23_n_87, ZN => L2_shift_L23_n_99);
  L2_shift_L23_g10696 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_77, A2 => L2_shift_L23_n_67, ZN => L2_shift_L23_n_98);
  L2_shift_L23_g10697 : ND2D1BWP7T port map(A1 => L2_shift_L23_n_76, A2 => L2_shift_L23_n_70, ZN => L2_shift_L23_n_97);
  L2_shift_L23_g10698 : INR2XD0BWP7T port map(A1 => L2_shift_L23_n_390, B1 => L2_shift_L23_n_394, ZN => L2_shift_gr_pos_load);
  L2_shift_L23_g10699 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_309, A2 => L2_shift_L23_n_312, A3 => L2_shift_L23_n_311, A4 => L2_shift_L23_n_310, ZN => L2_shift_L23_n_96);
  L2_shift_L23_g10700 : NR2D0BWP7T port map(A1 => L2_shift_L23_n_62, A2 => L2_shift_L23_n_84, ZN => L2_shift_L23_n_95);
  L2_shift_L23_g10701 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_396, A2 => L2_shift_L23_n_331, A3 => L2_shift_L23_n_290, A4 => L2_shift_L23_n_397, ZN => L2_shift_L23_n_94);
  L2_shift_L23_g10702 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_304, A2 => L2_shift_L23_n_308, A3 => L2_shift_L23_n_306, A4 => L2_shift_L23_n_307, ZN => L2_shift_L23_n_93);
  L2_shift_L23_g10703 : AOI221D0BWP7T port map(A1 => L2_shift_L23_n_309, A2 => L2_shift_L23_n_296, B1 => L2_shift_L23_n_310, B2 => L2_shift_L23_n_297, C => L2_shift_L23_n_79, ZN => L2_shift_L23_n_92);
  L2_shift_L23_g10704 : OR4D1BWP7T port map(A1 => L2_shift_L23_n_318, A2 => L2_shift_L23_n_320, A3 => L2_shift_L23_n_319, A4 => L2_shift_L23_n_317, Z => L2_shift_L23_n_91);
  L2_shift_L23_g10705 : AOI222D0BWP7T port map(A1 => L2_shift_L23_n_304, A2 => L2_shift_L23_n_60, B1 => L2_shift_L23_n_308, B2 => L2_shift_L23_n_296, C1 => L2_shift_L23_n_305, C2 => L2_shift_L23_n_58, ZN => L2_shift_L23_n_90);
  L2_shift_L23_g10706 : AOI222D0BWP7T port map(A1 => L2_shift_L23_n_315, A2 => L2_shift_L23_n_52, B1 => L2_shift_L23_n_314, B2 => L2_shift_L23_n_59, C1 => L2_shift_L23_n_313, C2 => L2_shift_L23_n_60, ZN => L2_shift_L23_n_89);
  L2_shift_L23_g10707 : INVD1BWP7T port map(I => L2_shift_L23_n_86, ZN => L2_shift_L23_n_85);
  L2_shift_L23_g10708 : NR3D0BWP7T port map(A1 => L2_shift_L23_n_313, A2 => L2_shift_L23_n_314, A3 => L2_shift_L23_n_315, ZN => L2_shift_L23_n_84);
  L2_shift_L23_g10709 : OR3D1BWP7T port map(A1 => L2_shift_L23_n_327, A2 => L2_shift_L23_n_328, A3 => L2_shift_L23_n_329, Z => L2_shift_L23_n_83);
  L2_shift_L23_g10710 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_323, A2 => L2_shift_L23_n_324, B => L2_shift_L23_n_61, ZN => L2_shift_L23_n_82);
  L2_shift_L23_g10711 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_303, A2 => L2_shift_L23_n_302, B => L2_shift_L23_n_292, ZN => L2_shift_L23_n_81);
  L2_shift_L23_g10712 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_52, A2 => L2_shift_L23_n_302, B1 => L2_shift_L23_n_303, B2 => L2_shift_L23_n_59, ZN => L2_shift_L23_n_80);
  L2_shift_L23_g10713 : AO22D0BWP7T port map(A1 => L2_shift_L23_n_312, A2 => L2_shift_L23_n_58, B1 => L2_shift_L23_n_282, B2 => L2_shift_L23_n_311, Z => L2_shift_L23_n_79);
  L2_shift_L23_g10714 : IND3D1BWP7T port map(A1 => cell_type_int(2), B1 => cell_type_int(1), B2 => L2_shift_L23_n_53, ZN => L2_shift_L23_n_394);
  L2_shift_L23_g10715 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_320, B1 => L2_shift_L23_n_397, B2 => L2_shift_L23_n_325, ZN => L2_shift_L23_n_88);
  L2_shift_L23_g10716 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_319, B1 => L2_shift_L23_n_397, B2 => L2_shift_L23_n_326, ZN => L2_shift_L23_n_87);
  L2_shift_L23_g10717 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_321, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_324, ZN => L2_shift_L23_n_86);
  L2_shift_L23_g10718 : INVD0BWP7T port map(I => L2_shift_L23_n_74, ZN => L2_shift_L23_n_73);
  L2_shift_L23_g10719 : INVD1BWP7T port map(I => L2_shift_L23_n_72, ZN => L2_shift_L23_n_71);
  L2_shift_L23_g10720 : INVD1BWP7T port map(I => L2_shift_L23_n_70, ZN => L2_shift_L23_n_69);
  L2_shift_L23_g10721 : INVD1BWP7T port map(I => L2_shift_L23_n_67, ZN => L2_shift_L23_n_68);
  L2_shift_L23_g10722 : INVD1BWP7T port map(I => L2_shift_L23_n_66, ZN => L2_shift_L23_n_65);
  L2_shift_L23_g10723 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_306, A2 => L2_shift_L23_n_282, B1 => L2_shift_L23_n_307, B2 => L2_shift_L23_n_297, ZN => L2_shift_L23_n_64);
  L2_shift_L23_g10724 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_289, A2 => L2_shift_L23_n_285, A3 => L2_shift_L23_n_283, A4 => L2_shift_L23_n_284, ZN => L2_shift_L23_n_63);
  L2_shift_L23_g10725 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_321, B1 => L2_shift_L23_n_397, B2 => L2_shift_L23_n_324, ZN => L2_shift_L23_n_78);
  L2_shift_L23_g10726 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_317, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_328, ZN => L2_shift_L23_n_77);
  L2_shift_L23_g10727 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_318, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_327, ZN => L2_shift_L23_n_76);
  L2_shift_L23_g10728 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_319, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_326, ZN => L2_shift_L23_n_75);
  L2_shift_L23_g10729 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_318, B1 => L2_shift_L23_n_397, B2 => L2_shift_L23_n_327, ZN => L2_shift_L23_n_74);
  L2_shift_L23_g10730 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_320, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_325, ZN => L2_shift_L23_n_72);
  L2_shift_L23_g10731 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_317, B1 => L2_shift_L23_n_397, B2 => L2_shift_L23_n_328, ZN => L2_shift_L23_n_70);
  L2_shift_L23_g10732 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_316, B1 => L2_shift_L23_n_397, B2 => L2_shift_L23_n_329, ZN => L2_shift_L23_n_67);
  L2_shift_L23_g10733 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_290, A2 => L2_shift_L23_n_322, B1 => L2_shift_L23_n_301, B2 => L2_shift_L23_n_323, ZN => L2_shift_L23_n_66);
  L2_shift_L23_g10734 : OR2D1BWP7T port map(A1 => L2_shift_L23_n_396, A2 => L2_shift_L23_n_301, Z => L2_shift_L23_n_62);
  L2_shift_L23_g10735 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_301, A2 => L2_shift_L23_n_397, ZN => L2_shift_L23_n_61);
  L2_shift_L23_g10736 : INVD0BWP7T port map(I => L2_shift_L23_n_298, ZN => L2_shift_L23_n_60);
  L2_shift_L23_g10738 : INVD0BWP7T port map(I => L2_county(2), ZN => L2_shift_L23_n_58);
  L2_shift_L23_g10739 : INVD1BWP7T port map(I => L2_pixel_array_to_shift(6), ZN => L2_shift_L23_n_57);
  L2_shift_L23_g10740 : INVD1BWP7T port map(I => L2_pixel_array_to_shift(1), ZN => L2_shift_L23_n_56);
  L2_shift_L23_g10741 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(2), ZN => L2_shift_L23_n_55);
  L2_shift_L23_g10742 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(3), ZN => L2_shift_L23_n_54);
  L2_shift_L23_g10743 : CKND1BWP7T port map(I => cell_type_int(0), ZN => L2_shift_L23_n_53);
  L2_shift_L23_g10744 : INVD0BWP7T port map(I => L2_shift_L23_n_300, ZN => L2_shift_L23_n_52);
  L2_shift_L23_g10745 : CKND1BWP7T port map(I => L2_pixel_array_to_shift(7), ZN => L2_shift_L23_n_51);
  L2_shift_L23_g10746 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(4), ZN => L2_shift_L23_n_50);
  L2_shift_L23_g10747 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(5), ZN => L2_shift_L23_n_49);
  L2_shift_L23_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L23_n_48, Q => L2_shift_L23_state(0));
  L2_shift_L23_g10066 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_47, A2 => L2_shift_L23_n_6, A3 => L2_shift_L23_n_15, A4 => reset, ZN => L2_shift_L23_n_48);
  L2_shift_L23_g10068 : OAI211D1BWP7T port map(A1 => L2_shift_L23_n_2, A2 => L2_shift_L23_n_5, B => L2_shift_L23_n_18, C => L2_shift_L23_n_45, ZN => L2_shift_L23_n_47);
  L2_shift_L23_g10069 : ND4D0BWP7T port map(A1 => L2_shift_L23_n_26, A2 => L2_shift_L23_n_25, A3 => L2_shift_L23_n_41, A4 => L2_shift_L23_n_27, ZN => L2_shift_L23_n_46);
  L2_shift_L23_g10070 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_42, A2 => L2_shift_shift_pulse_gr, B1 => L2_shift_L23_n_32, B2 => L2_shift_shift_pulse_gr, ZN => L2_shift_L23_n_45);
  L2_shift_L23_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L23_n_44, Q => L2_shift_L23_state(1));
  L2_shift_L23_g10073 : IND4D0BWP7T port map(A1 => L2_shift_L23_n_15, B1 => L2_shift_L23_n_13, B2 => L2_shift_L23_n_26, B3 => L2_shift_L23_n_39, ZN => L2_shift_L23_n_44);
  L2_shift_L23_g10074 : IND4D0BWP7T port map(A1 => L2_shift_L23_n_38, B1 => L2_shift_L23_n_17, B2 => L2_shift_L23_n_13, B3 => L2_shift_L23_n_16, ZN => L2_shift_L23_n_43);
  L2_shift_L23_g10075 : IINR4D0BWP7T port map(A1 => L2_shift_L23_n_37, A2 => L2_shift_L23_n_5, B1 => L2_shift_L23_n_390, B2 => L2_shift_L23_n_316, ZN => L2_shift_L23_n_42);
  L2_shift_L23_state_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L23_n_40, Q => L2_shift_L23_state(2));
  L2_shift_L23_g10077 : AOI221D0BWP7T port map(A1 => L2_shift_L23_n_36, A2 => L2_shift_L23_n_1, B1 => L2_shift_L23_n_316, B2 => L2_shift_L23_n_4, C => L2_shift_L23_n_20, ZN => L2_shift_L23_n_41);
  L2_shift_L23_g10078 : IND4D0BWP7T port map(A1 => L2_shift_L23_n_29, B1 => L2_shift_L23_n_27, B2 => L2_shift_L23_n_31, B3 => L2_shift_L23_n_33, ZN => L2_shift_L23_n_40);
  L2_shift_L23_g10079 : NR3D0BWP7T port map(A1 => L2_shift_L23_n_24, A2 => L2_shift_L23_n_34, A3 => L2_shift_L23_n_29, ZN => L2_shift_L23_n_39);
  L2_shift_L23_g10080 : ND4D0BWP7T port map(A1 => L2_shift_L23_n_30, A2 => L2_shift_L23_n_25, A3 => L2_shift_L23_n_31, A4 => L2_shift_L23_n_19, ZN => L2_shift_L23_n_38);
  L2_shift_L23_g10081 : INR4D0BWP7T port map(A1 => L2_shift_L23_n_32, B1 => L2_shift_L23_n_302, B2 => L2_shift_L23_n_330, B3 => L2_shift_gr_pos_reset, ZN => L2_shift_L23_n_37);
  L2_shift_L23_g10082 : IND2D1BWP7T port map(A1 => L2_shift_L23_n_328, B1 => L2_shift_L23_n_35, ZN => L2_shift_L23_n_36);
  L2_shift_L23_g10083 : NR4D0BWP7T port map(A1 => L2_shift_L23_n_22, A2 => L2_shift_L23_n_312, A3 => L2_shift_L23_n_314, A4 => L2_shift_L23_n_310, ZN => L2_shift_L23_n_35);
  L2_shift_L23_g10084 : AO221D0BWP7T port map(A1 => L2_shift_L23_n_28, A2 => L2_shift_shift_pulse_gr, B1 => L2_shift_L23_n_23, B2 => L2_shift_L23_n_2, C => L2_shift_L23_n_21, Z => L2_shift_L23_n_34);
  L2_shift_L23_g10085 : AOI222D0BWP7T port map(A1 => L2_shift_L23_n_23, A2 => L2_shift_shift_pulse_gr, B1 => L2_shift_L23_n_7, B2 => L2_shift_L23_n_1, C1 => L2_shift_L23_n_318, C2 => L2_shift_L23_n_4, ZN => L2_shift_L23_n_33);
  L2_shift_L23_g10086 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_28, A2 => L2_shift_L23_n_23, ZN => L2_shift_L23_n_32);
  L2_shift_L23_g10087 : AOI222D0BWP7T port map(A1 => L2_shift_L23_n_11, A2 => L2_shift_L23_n_396, B1 => L2_shift_L23_n_323, B2 => L2_shift_L23_n_4, C1 => L2_shift_L23_n_8, C2 => L2_shift_L23_n_1, ZN => L2_shift_L23_n_30);
  L2_shift_L23_g10088 : AOI211XD0BWP7T port map(A1 => L2_shift_L23_n_305, A2 => L2_shift_L23_n_1, B => L2_shift_L23_n_12, C => L2_shift_L23_n_20, ZN => L2_shift_L23_n_31);
  L2_shift_L23_g10089 : IOA21D1BWP7T port map(A1 => L2_shift_L23_n_319, A2 => L2_shift_L23_n_1, B => L2_shift_L23_n_19, ZN => L2_shift_L23_n_29);
  L2_shift_L23_g10090 : IND3D1BWP7T port map(A1 => L2_shift_L23_n_12, B1 => L2_shift_L23_n_10, B2 => L2_shift_L23_n_17, ZN => L2_shift_L23_n_28);
  L2_shift_L23_g10091 : MAOI22D0BWP7T port map(A1 => L2_shift_L23_n_324, A2 => L2_shift_L23_n_4, B1 => L2_shift_L23_n_14, B2 => reset, ZN => L2_shift_L23_n_27);
  L2_shift_L23_g10092 : MOAI22D0BWP7T port map(A1 => L2_shift_L23_n_5, A2 => L2_shift_L23_n_3, B1 => L2_shift_L23_n_11, B2 => L2_shift_L23_n_397, ZN => L2_shift_L23_n_24);
  L2_shift_L23_g10093 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_11, A2 => L2_shift_L23_n_290, B1 => L2_shift_L23_n_329, B2 => L2_shift_L23_n_1, ZN => L2_shift_L23_n_26);
  L2_shift_L23_g10094 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_11, A2 => L2_shift_L23_n_331, B1 => L2_shift_L23_n_315, B2 => L2_shift_L23_n_1, ZN => L2_shift_L23_n_25);
  L2_shift_L23_g10095 : AO211D0BWP7T port map(A1 => L2_shift_L23_n_318, A2 => L2_shift_shift_pulse_gr, B => L2_shift_L23_n_313, C => L2_shift_L23_n_317, Z => L2_shift_L23_n_22);
  L2_shift_L23_g10096 : OA21D0BWP7T port map(A1 => L2_shift_L23_n_6, A2 => L2_shift_L23_n_325, B => L2_shift_L23_n_1, Z => L2_shift_L23_n_21);
  L2_shift_L23_g10097 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_9, A2 => reset, B => L2_shift_L23_n_16, ZN => L2_shift_L23_n_23);
  L2_shift_L23_g10098 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_331, A2 => L2_shift_L23_n_290, B => L2_shift_L23_n_11, ZN => L2_shift_L23_n_18);
  L2_shift_L23_g10099 : AO21D0BWP7T port map(A1 => L2_shift_L23_n_311, A2 => L2_shift_L23_n_1, B => L2_shift_L23_n_15, Z => L2_shift_L23_n_20);
  L2_shift_L23_g10100 : AOI22D0BWP7T port map(A1 => L2_shift_L23_n_302, A2 => L2_shift_L23_n_4, B1 => L2_shift_L23_n_303, B2 => L2_shift_L23_n_1, ZN => L2_shift_L23_n_19);
  L2_shift_L23_g10101 : NR3D0BWP7T port map(A1 => L2_shift_L23_n_325, A2 => L2_shift_L23_n_326, A3 => L2_shift_L23_n_327, ZN => L2_shift_L23_n_14);
  L2_shift_L23_g10102 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_314, A2 => L2_shift_L23_n_308, B => L2_shift_L23_n_1, ZN => L2_shift_L23_n_17);
  L2_shift_L23_g10103 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_312, A2 => L2_shift_L23_n_306, B => L2_shift_L23_n_1, ZN => L2_shift_L23_n_16);
  L2_shift_L23_g10104 : AN2D1BWP7T port map(A1 => L2_shift_L23_n_309, A2 => L2_shift_L23_n_4, Z => L2_shift_L23_n_15);
  L2_shift_L23_g10105 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_320, A2 => L2_shift_L23_n_326, B => L2_shift_L23_n_1, ZN => L2_shift_L23_n_10);
  L2_shift_L23_g10106 : OAI21D0BWP7T port map(A1 => L2_shift_L23_n_313, A2 => L2_shift_L23_n_307, B => L2_shift_L23_n_1, ZN => L2_shift_L23_n_13);
  L2_shift_L23_g10107 : OA21D0BWP7T port map(A1 => L2_shift_L23_n_304, A2 => L2_shift_L23_n_310, B => L2_shift_L23_n_1, Z => L2_shift_L23_n_12);
  L2_shift_L23_g10108 : INR3D0BWP7T port map(A1 => L2_shift_L23_n_390, B1 => reset, B2 => L2_shift_L23_n_394, ZN => L2_shift_L23_n_11);
  L2_shift_L23_g10109 : NR2D0BWP7T port map(A1 => L2_shift_L23_n_328, A2 => L2_shift_L23_n_322, ZN => L2_shift_L23_n_9);
  L2_shift_L23_g10110 : AN2D0BWP7T port map(A1 => L2_shift_L23_n_324, A2 => L2_shift_shift_pulse_gr, Z => L2_shift_L23_n_8);
  L2_shift_L23_g10111 : OR2D1BWP7T port map(A1 => L2_shift_L23_n_320, A2 => L2_shift_L23_n_321, Z => L2_shift_L23_n_7);
  L2_shift_L23_g10112 : INVD0BWP7T port map(I => L2_shift_L23_n_4, ZN => L2_shift_L23_n_3);
  L2_shift_L23_g10113 : INR2D1BWP7T port map(A1 => L2_shift_L23_n_330, B1 => L2_calc_start_internal, ZN => L2_shift_L23_n_6);
  L2_shift_L23_g10114 : NR2D1BWP7T port map(A1 => L2_shift_L23_n_318, A2 => L2_shift_L23_n_324, ZN => L2_shift_L23_n_5);
  L2_shift_L23_g10115 : NR2D1BWP7T port map(A1 => reset, A2 => L2_shift_shift_pulse_gr, ZN => L2_shift_L23_n_4);
  L2_shift_L23_g10116 : INVD0BWP7T port map(I => L2_shift_shift_pulse_gr, ZN => L2_shift_L23_n_2);
  L2_shift_L23_drc_bufs10119 : INVD0BWP7T port map(I => reset, ZN => L2_shift_L23_n_1);
  L2_shift_L23_state_reg_3 : DFD1BWP7T port map(CP => clk, D => L2_shift_L23_n_46, Q => L2_shift_L23_state(3), QN => L2_shift_L23_n_146);
  L2_shift_L23_state_reg_4 : DFD1BWP7T port map(CP => clk, D => L2_shift_L23_n_43, Q => L2_shift_L23_state(4), QN => L2_shift_L23_n_145);
  L2_shift_L23_g17815 : INR4D0BWP7T port map(A1 => L2_shift_L23_n_253, B1 => L2_shift_L23_n_129, B2 => L2_shift_L23_n_288, B3 => L2_shift_L23_n_110, ZN => L2_shift_L23_n_398);
  L2_shift_L23_g17816 : OA222D0BWP7T port map(A1 => L2_shift_L23_n_262, A2 => L2_shift_L23_n_182, B1 => L2_shift_L23_n_259, B2 => L2_shift_L23_n_208, C1 => L2_shift_L23_n_256, C2 => L2_shift_L23_n_181, Z => L2_shift_L23_n_399);
  L2_gameovercontrol_go_type_reg_0 : DFKSND1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_123, SN => L2_gameovercontrol_n_93, Q => L2_in_go_sprite_type(0), QN => UNCONNECTED2);
  L2_gameovercontrol_go_type_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_129, Q => L2_in_go_sprite_type(1));
  L2_gameovercontrol_go_type_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_127, Q => L2_in_go_sprite_type(2));
  L2_gameovercontrol_go_type_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_126, Q => L2_in_go_sprite_type(3));
  L2_gameovercontrol_go_type_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_122, Q => L2_in_go_sprite_type(4));
  L2_gameovercontrol_g4073 : IND4D0BWP7T port map(A1 => L2_gameovercontrol_n_128, B1 => L2_gameovercontrol_n_118, B2 => L2_gameovercontrol_n_117, B3 => L2_gameovercontrol_n_116, ZN => L2_gameovercontrol_n_129);
  L2_gameovercontrol_g4075 : OAI211D1BWP7T port map(A1 => L2_current_block_horizontal(1), A2 => L2_gameovercontrol_n_111, B => L2_gameovercontrol_n_125, C => L2_gameovercontrol_n_96, ZN => L2_gameovercontrol_n_128);
  L2_gameovercontrol_g4076 : ND3D0BWP7T port map(A1 => L2_gameovercontrol_n_124, A2 => L2_gameovercontrol_n_115, A3 => L2_gameovercontrol_n_66, ZN => L2_gameovercontrol_n_127);
  L2_gameovercontrol_g4080 : IND4D0BWP7T port map(A1 => L2_gameovercontrol_n_120, B1 => L2_gameovercontrol_n_109, B2 => L2_gameovercontrol_n_106, B3 => L2_gameovercontrol_n_118, ZN => L2_gameovercontrol_n_126);
  L2_gameovercontrol_g4081 : AOI31D0BWP7T port map(A1 => L2_gameovercontrol_n_100, A2 => L2_gameovercontrol_n_46, A3 => L2_in_score_12bits(9), B => L2_gameovercontrol_n_121, ZN => L2_gameovercontrol_n_125);
  L2_gameovercontrol_g4082 : AOI221D0BWP7T port map(A1 => L2_gameovercontrol_n_113, A2 => L2_in_st_go_sel, B1 => L2_gameovercontrol_n_80, B2 => L2_gameovercontrol_n_46, C => L2_gameovercontrol_n_103, ZN => L2_gameovercontrol_n_124);
  L2_gameovercontrol_g4083 : AN2D1BWP7T port map(A1 => L2_in_go_colour(2), A2 => L2_gameovercontrol_n_55, Z => L2_in_go_colour(1));
  L2_gameovercontrol_g4084 : OAI211D1BWP7T port map(A1 => reset, A2 => L2_gameovercontrol_n_91, B => L2_gameovercontrol_n_112, C => L2_gameovercontrol_n_102, ZN => L2_gameovercontrol_n_123);
  L2_gameovercontrol_g4085 : OAI221D0BWP7T port map(A1 => L2_gameovercontrol_n_89, A2 => L2_gameovercontrol_n_62, B1 => L2_gameovercontrol_row, B2 => L2_gameovercontrol_n_107, C => L2_gameovercontrol_n_93, ZN => L2_gameovercontrol_n_122);
  L2_gameovercontrol_g4086 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_119, A2 => L2_gameovercontrol_n_54, B => L2_gameovercontrol_n_131, ZN => L2_reset_county_go);
  L2_gameovercontrol_g4087 : OAI22D0BWP7T port map(A1 => L2_gameovercontrol_n_114, A2 => L2_current_block_horizontal(0), B1 => L2_gameovercontrol_n_99, B2 => L2_current_block_horizontal(1), ZN => L2_gameovercontrol_n_121);
  L2_gameovercontrol_g4088 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_119, A2 => L2_gameovercontrol_n_164, ZN => L2_gameovercontrol_n_162);
  L2_gameovercontrol_g4089 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_110, A2 => L2_gameovercontrol_n_54, B => L2_gameovercontrol_n_131, ZN => L2_reset_dual_pixel_y_go);
  L2_gameovercontrol_g4090 : NR3D0BWP7T port map(A1 => L2_gameovercontrol_n_110, A2 => L2_gameovercontrol_n_164, A3 => L2_gameovercontrol_n_71, ZN => L2_en_county_go);
  L2_gameovercontrol_g4091 : OAI222D0BWP7T port map(A1 => L2_gameovercontrol_n_92, A2 => L2_gameovercontrol_n_76, B1 => L2_gameovercontrol_n_58, B2 => L2_gameovercontrol_n_111, C1 => L2_gameovercontrol_row, C2 => L2_gameovercontrol_n_101, ZN => L2_gameovercontrol_n_120);
  L2_gameovercontrol_g4092 : OAI22D0BWP7T port map(A1 => L2_gameovercontrol_n_104, A2 => L2_gameovercontrol_state(0), B1 => L2_gameovercontrol_n_90, B2 => L2_gameovercontrol_n_65, ZN => L2_in_go_colour(2));
  L2_gameovercontrol_g4093 : OAI211D1BWP7T port map(A1 => L2_in_score_12bits(1), A2 => L2_gameovercontrol_n_42, B => L2_gameovercontrol_n_100, C => L2_gameovercontrol_n_60, ZN => L2_gameovercontrol_n_117);
  L2_gameovercontrol_g4094 : IND3D1BWP7T port map(A1 => L2_gameovercontrol_n_99, B1 => L2_in_score_12bits(5), B2 => L2_current_block_horizontal(2), ZN => L2_gameovercontrol_n_116);
  L2_gameovercontrol_g4095 : NR3D0BWP7T port map(A1 => L2_gameovercontrol_n_165, A2 => L2_gameovercontrol_n_164, A3 => L2_dual_pixel_y, ZN => L2_en_dual_pixel_y_go);
  L2_gameovercontrol_g4096 : IND2D1BWP7T port map(A1 => L2_gameovercontrol_n_110, B1 => L2_gameovercontrol_n_71, ZN => L2_gameovercontrol_n_119);
  L2_gameovercontrol_g4097 : ND3D0BWP7T port map(A1 => L2_gameovercontrol_n_95, A2 => L2_in_st_go_sel, A3 => L2_gameovercontrol_row, ZN => L2_gameovercontrol_n_118);
  L2_gameovercontrol_g4098 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_165, A2 => L2_gameovercontrol_n_54, B => L2_gameovercontrol_n_131, ZN => L2_reset_current_block_horizontal_go);
  L2_gameovercontrol_g4099 : AOI21D0BWP7T port map(A1 => L2_gameovercontrol_n_64, A2 => L2_gameovercontrol_n_59, B => L2_gameovercontrol_n_108, ZN => L2_gameovercontrol_n_115);
  L2_gameovercontrol_g4100 : OA21D0BWP7T port map(A1 => L2_gameovercontrol_n_97, A2 => L2_gameovercontrol_row, B => L2_gameovercontrol_n_101, Z => L2_gameovercontrol_n_114);
  L2_gameovercontrol_g4101 : OAI22D0BWP7T port map(A1 => L2_gameovercontrol_n_94, A2 => reset, B1 => L2_gameovercontrol_n_75, B2 => L2_gameovercontrol_n_48, ZN => L2_gameovercontrol_n_113);
  L2_gameovercontrol_g4102 : AOI31D0BWP7T port map(A1 => L2_gameovercontrol_n_56, A2 => L2_gameovercontrol_n_60, A3 => L2_gameovercontrol_n_47, B => L2_gameovercontrol_n_105, ZN => L2_gameovercontrol_n_112);
  L2_gameovercontrol_g4103 : IOA21D0BWP7T port map(A1 => L2_gameovercontrol_n_82, A2 => L2_gameovercontrol_n_53, B => L2_gameovercontrol_n_100, ZN => L2_gameovercontrol_n_109);
  L2_gameovercontrol_g4104 : INR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_165, B1 => L2_gameovercontrol_n_164, ZN => L2_en_current_block_horizontal_go);
  L2_gameovercontrol_g4105 : AOI31D0BWP7T port map(A1 => L2_gameovercontrol_n_73, A2 => L2_gameovercontrol_n_49, A3 => L2_current_block_horizontal(3), B => L2_gameovercontrol_n_62, ZN => L2_gameovercontrol_n_108);
  L2_gameovercontrol_g4106 : ND3D0BWP7T port map(A1 => L2_gameovercontrol_n_87, A2 => L2_current_block_horizontal(0), A3 => L2_gameovercontrol_row, ZN => L2_gameovercontrol_n_111);
  L2_gameovercontrol_g4107 : IND2D1BWP7T port map(A1 => L2_gameovercontrol_n_165, B1 => L2_dual_pixel_y, ZN => L2_gameovercontrol_n_110);
  L2_gameovercontrol_g4108 : IAO21D0BWP7T port map(A1 => L2_gameovercontrol_n_84, A2 => reset, B => L2_gameovercontrol_n_64, ZN => L2_gameovercontrol_n_107);
  L2_gameovercontrol_g4109 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_42, A2 => L2_in_score_12bits(7), B => L2_gameovercontrol_n_98, ZN => L2_gameovercontrol_n_106);
  L2_gameovercontrol_g4110 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_81, A2 => L2_gameovercontrol_n_62, B => L2_gameovercontrol_n_85, ZN => L2_gameovercontrol_n_105);
  L2_gameovercontrol_g4111 : AOI22D0BWP7T port map(A1 => L2_gameovercontrol_n_83, A2 => L2_gameovercontrol_state(2), B1 => L2_gameovercontrol_n_79, B2 => L2_gameovercontrol_pixel_arr_buffer(6), ZN => L2_gameovercontrol_n_104);
  L2_gameovercontrol_g4112 : AO33D0BWP7T port map(A1 => L2_gameovercontrol_n_56, A2 => L2_gameovercontrol_n_68, A3 => L2_gameovercontrol_n_47, B1 => L2_gameovercontrol_n_80, B2 => L2_current_block_horizontal(2), B3 => L2_in_score_12bits(6), Z => L2_gameovercontrol_n_103);
  L2_gameovercontrol_g4113 : AOI32D1BWP7T port map(A1 => L2_gameovercontrol_n_78, A2 => L2_gameovercontrol_n_47, A3 => L2_in_score_12bits(0), B1 => L2_gameovercontrol_n_74, B2 => L2_gameovercontrol_n_61, ZN => L2_gameovercontrol_n_102);
  L2_gameovercontrol_g4114 : CKND1BWP7T port map(I => L2_gameovercontrol_n_98, ZN => L2_gameovercontrol_n_99);
  L2_gameovercontrol_g4115 : AOI21D0BWP7T port map(A1 => L2_gameovercontrol_n_77, A2 => L2_current_block_horizontal(1), B => L2_gameovercontrol_n_87, ZN => L2_gameovercontrol_n_97);
  L2_gameovercontrol_g4116 : IND4D0BWP7T port map(A1 => L2_gameovercontrol_n_58, B1 => L2_current_block_horizontal(0), B2 => L2_gameovercontrol_n_77, B3 => L2_gameovercontrol_n_56, ZN => L2_gameovercontrol_n_96);
  L2_gameovercontrol_g4117 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_86, A2 => L2_current_block_horizontal(4), ZN => L2_gameovercontrol_n_95);
  L2_gameovercontrol_g4118 : AOI31D0BWP7T port map(A1 => L2_gameovercontrol_n_46, A2 => L2_gameovercontrol_row, A3 => L2_in_score_12bits(10), B => L2_gameovercontrol_n_52, ZN => L2_gameovercontrol_n_94);
  L2_gameovercontrol_g4119 : IND2D1BWP7T port map(A1 => L2_gameovercontrol_n_53, B1 => L2_gameovercontrol_n_87, ZN => L2_gameovercontrol_n_101);
  L2_gameovercontrol_g4120 : NR2D1BWP7T port map(A1 => L2_gameovercontrol_n_88, A2 => L2_gameovercontrol_n_40, ZN => L2_gameovercontrol_n_100);
  L2_gameovercontrol_g4121 : NR2D1BWP7T port map(A1 => L2_gameovercontrol_n_88, A2 => L2_gameovercontrol_n_51, ZN => L2_gameovercontrol_n_98);
  L2_gameovercontrol_g4122 : AOI22D0BWP7T port map(A1 => L2_gameovercontrol_n_56, A2 => L2_gameovercontrol_n_74, B1 => L2_gameovercontrol_n_50, B2 => L2_gameovercontrol_n_46, ZN => L2_gameovercontrol_n_92);
  L2_gameovercontrol_g4123 : AOI32D1BWP7T port map(A1 => L2_gameovercontrol_n_46, A2 => L2_gameovercontrol_row, A3 => L2_in_score_12bits(8), B1 => L2_gameovercontrol_n_72, B2 => L2_in_st_go_sel, ZN => L2_gameovercontrol_n_91);
  L2_gameovercontrol_g4124 : AOI32D1BWP7T port map(A1 => L2_gameovercontrol_n_3, A2 => L2_gameovercontrol_state(2), A3 => L2_gameovercontrol_pixel_arr_buffer(3), B1 => L2_gameovercontrol_n_67, B2 => L2_gameovercontrol_state(1), ZN => L2_gameovercontrol_n_90);
  L2_gameovercontrol_g4125 : AOI222D0BWP7T port map(A1 => L2_gameovercontrol_n_50, A2 => L2_gameovercontrol_n_42, B1 => L2_gameovercontrol_n_51, B2 => L2_current_block_horizontal(2), C1 => L2_gameovercontrol_row, C2 => L2_current_block_horizontal(1), ZN => L2_gameovercontrol_n_89);
  L2_gameovercontrol_g4126 : OA21D0BWP7T port map(A1 => L2_gameovercontrol_n_78, A2 => L2_gameovercontrol_n_63, B => L2_gameovercontrol_n_66, Z => L2_gameovercontrol_n_93);
  L2_gameovercontrol_g4127 : IND3D1BWP7T port map(A1 => L2_gameovercontrol_n_79, B1 => L2_gameovercontrol_n_65, B2 => L2_gameovercontrol_n_69, ZN => L2_gameovercontrol_n_131);
  L2_gameovercontrol_g4128 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_78, A2 => L2_current_block_horizontal(3), B => L2_current_block_horizontal(4), ZN => L2_gameovercontrol_n_165);
  L2_gameovercontrol_g4129 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_78, A2 => L2_gameovercontrol_n_64, ZN => L2_gameovercontrol_n_86);
  L2_gameovercontrol_g4130 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_77, A2 => L2_in_st_go_sel, ZN => L2_gameovercontrol_n_88);
  L2_gameovercontrol_g4131 : NR2D1BWP7T port map(A1 => L2_gameovercontrol_n_76, A2 => L2_in_st_go_sel, ZN => L2_gameovercontrol_n_87);
  L2_gameovercontrol_g4132 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_79, A2 => L2_gameovercontrol_state(0), ZN => L2_gameovercontrol_n_164);
  L2_gameovercontrol_g4133 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_49, A2 => L2_in_score_12bits(4), B => L2_gameovercontrol_n_80, ZN => L2_gameovercontrol_n_85);
  L2_gameovercontrol_g4134 : AOI21D0BWP7T port map(A1 => L2_gameovercontrol_n_49, A2 => L2_current_block_horizontal(0), B => L2_gameovercontrol_n_57, ZN => L2_gameovercontrol_n_84);
  L2_gameovercontrol_g4135 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_70, A2 => L2_gameovercontrol_state(3), ZN => L2_gameovercontrol_n_83);
  L2_gameovercontrol_g4136 : AOI22D0BWP7T port map(A1 => L2_gameovercontrol_n_46, A2 => L2_in_score_12bits(11), B1 => L2_gameovercontrol_n_60, B2 => L2_in_score_12bits(3), ZN => L2_gameovercontrol_n_82);
  L2_gameovercontrol_g4137 : AOI32D1BWP7T port map(A1 => L2_gameovercontrol_n_40, A2 => L2_gameovercontrol_n_41, A3 => L2_current_block_horizontal(0), B1 => L2_gameovercontrol_n_58, B2 => L2_gameovercontrol_row, ZN => L2_gameovercontrol_n_81);
  L2_gameovercontrol_g4138 : CKND1BWP7T port map(I => L2_gameovercontrol_n_77, ZN => L2_gameovercontrol_n_76);
  L2_gameovercontrol_g4139 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_60, A2 => L2_in_score_12bits(2), ZN => L2_gameovercontrol_n_75);
  L2_gameovercontrol_g4140 : OR2D1BWP7T port map(A1 => L2_gameovercontrol_n_65, A2 => L2_gameovercontrol_state(2), Z => L2_gameovercontrol_n_976_BAR);
  L2_gameovercontrol_g4141 : NR2D1BWP7T port map(A1 => L2_gameovercontrol_n_51, A2 => reset, ZN => L2_gameovercontrol_n_80);
  L2_gameovercontrol_g4142 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_163, A2 => L2_gameovercontrol_state(1), ZN => L2_gameovercontrol_n_79);
  L2_gameovercontrol_g4143 : NR2D1BWP7T port map(A1 => L2_gameovercontrol_n_49, A2 => L2_gameovercontrol_n_43, ZN => L2_gameovercontrol_n_78);
  L2_gameovercontrol_g4144 : NR2D1BWP7T port map(A1 => L2_gameovercontrol_n_48, A2 => L2_current_block_horizontal(4), ZN => L2_gameovercontrol_n_77);
  L2_gameovercontrol_g4145 : CKND1BWP7T port map(I => L2_gameovercontrol_n_72, ZN => L2_gameovercontrol_n_73);
  L2_gameovercontrol_g4146 : AOI22D0BWP7T port map(A1 => L2_gameovercontrol_n_3, A2 => L2_gameovercontrol_pixel_arr_buffer(2), B1 => L2_gameovercontrol_state(1), B2 => L2_gameovercontrol_pixel_arr_buffer(4), ZN => L2_gameovercontrol_n_70);
  L2_gameovercontrol_g4147 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_state(1), A2 => L2_gameovercontrol_state(2), B => L2_gameovercontrol_n_45, ZN => L2_gameovercontrol_n_69);
  L2_gameovercontrol_g4148 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_43, A2 => L2_gameovercontrol_n_42, B => L2_gameovercontrol_n_41, ZN => L2_gameovercontrol_n_68);
  L2_gameovercontrol_g4149 : MUX2D1BWP7T port map(I0 => L2_gameovercontrol_pixel_arr_buffer(1), I1 => L2_gameovercontrol_pixel_arr_buffer(5), S => L2_gameovercontrol_state(2), Z => L2_gameovercontrol_n_67);
  L2_gameovercontrol_g4150 : OAI21D0BWP7T port map(A1 => L2_gameovercontrol_n_41, A2 => L2_current_block_horizontal(0), B => L2_gameovercontrol_n_49, ZN => L2_gameovercontrol_n_74);
  L2_gameovercontrol_g4151 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_58, A2 => L2_current_block_horizontal(0), ZN => L2_gameovercontrol_n_72);
  L2_gameovercontrol_g4152 : AN3D1BWP7T port map(A1 => L2_county(0), A2 => L2_county(2), A3 => L2_in_go_y_pos(1), Z => L2_gameovercontrol_n_71);
  L2_gameovercontrol_g4153 : INVD0BWP7T port map(I => L2_gameovercontrol_n_64, ZN => L2_gameovercontrol_n_63);
  L2_gameovercontrol_g4154 : INVD0BWP7T port map(I => L2_gameovercontrol_n_61, ZN => L2_gameovercontrol_n_62);
  L2_gameovercontrol_g4155 : INVD0BWP7T port map(I => L2_gameovercontrol_n_60, ZN => L2_gameovercontrol_n_59);
  L2_gameovercontrol_g4156 : INVD0BWP7T port map(I => L2_gameovercontrol_n_58, ZN => L2_gameovercontrol_n_57);
  L2_gameovercontrol_g4157 : INVD1BWP7T port map(I => L2_gameovercontrol_n_55, ZN => L2_gameovercontrol_n_56);
  L2_gameovercontrol_g4158 : IND2D1BWP7T port map(A1 => reset, B1 => L2_current_block_horizontal(4), ZN => L2_gameovercontrol_n_66);
  L2_gameovercontrol_g4159 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_45, A2 => L2_gameovercontrol_state(0), ZN => L2_gameovercontrol_n_65);
  L2_gameovercontrol_g4160 : NR2XD0BWP7T port map(A1 => L2_current_block_horizontal(3), A2 => reset, ZN => L2_gameovercontrol_n_64);
  L2_gameovercontrol_g4161 : NR2D1BWP7T port map(A1 => L2_in_st_go_sel, A2 => reset, ZN => L2_gameovercontrol_n_61);
  L2_gameovercontrol_g4162 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_41, A2 => L2_gameovercontrol_n_43, ZN => L2_gameovercontrol_n_60);
  L2_gameovercontrol_g4163 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_41, A2 => L2_gameovercontrol_n_42, ZN => L2_gameovercontrol_n_58);
  L2_gameovercontrol_g4164 : ND2D1BWP7T port map(A1 => L2_in_st_go_sel, A2 => L2_gameovercontrol_n_40, ZN => L2_gameovercontrol_n_55);
  L2_gameovercontrol_g4165 : INVD0BWP7T port map(I => L2_gameovercontrol_n_53, ZN => L2_gameovercontrol_n_52);
  L2_gameovercontrol_g4166 : INVD0BWP7T port map(I => L2_gameovercontrol_n_51, ZN => L2_gameovercontrol_n_50);
  L2_gameovercontrol_g4167 : INVD0BWP7T port map(I => L2_gameovercontrol_n_48, ZN => L2_gameovercontrol_n_47);
  L2_gameovercontrol_g4168 : IND2D1BWP7T port map(A1 => L2_gameovercontrol_state(2), B1 => L2_gameovercontrol_state(3), ZN => L2_gameovercontrol_n_163);
  L2_gameovercontrol_g4169 : CKND2D1BWP7T port map(A1 => L2_gameovercontrol_state(0), A2 => L2_gameovercontrol_state(3), ZN => L2_gameovercontrol_n_54);
  L2_gameovercontrol_g4170 : CKND2D1BWP7T port map(A1 => L2_gameovercontrol_n_42, A2 => L2_current_block_horizontal(1), ZN => L2_gameovercontrol_n_53);
  L2_gameovercontrol_g4171 : CKND2D1BWP7T port map(A1 => L2_gameovercontrol_n_43, A2 => L2_gameovercontrol_row, ZN => L2_gameovercontrol_n_51);
  L2_gameovercontrol_g4172 : CKND2D1BWP7T port map(A1 => L2_current_block_horizontal(2), A2 => L2_current_block_horizontal(1), ZN => L2_gameovercontrol_n_49);
  L2_gameovercontrol_g4173 : IND2D1BWP7T port map(A1 => reset, B1 => L2_current_block_horizontal(3), ZN => L2_gameovercontrol_n_48);
  L2_gameovercontrol_g4174 : NR2D1BWP7T port map(A1 => L2_gameovercontrol_n_42, A2 => L2_current_block_horizontal(1), ZN => L2_gameovercontrol_n_46);
  L2_gameovercontrol_g4177 : INVD1BWP7T port map(I => L2_current_block_horizontal(0), ZN => L2_gameovercontrol_n_43);
  L2_gameovercontrol_g4178 : INVD1BWP7T port map(I => L2_current_block_horizontal(2), ZN => L2_gameovercontrol_n_42);
  L2_gameovercontrol_g4179 : INVD1BWP7T port map(I => L2_current_block_horizontal(1), ZN => L2_gameovercontrol_n_41);
  L2_gameovercontrol_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_37, Q => L2_gameovercontrol_state(0));
  L2_gameovercontrol_g3220 : AO211D0BWP7T port map(A1 => L2_gameovercontrol_n_22, A2 => L2_gameovercontrol_n_9, B => L2_gameovercontrol_n_166, C => L2_gameovercontrol_n_31, Z => L2_gameovercontrol_n_37);
  L2_gameovercontrol_g3221 : IOA21D1BWP7T port map(A1 => L2_gameovercontrol_n_31, A2 => L2_gameovercontrol_state(1), B => L2_gameovercontrol_n_34, ZN => L2_gameovercontrol_n_36);
  L2_gameovercontrol_state_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_32, Q => L2_gameovercontrol_state(2));
  L2_gameovercontrol_g3223 : AO21D0BWP7T port map(A1 => L2_gameovercontrol_n_27, A2 => L2_gameovercontrol_n_6, B => L2_gameovercontrol_n_166, Z => L2_gameovercontrol_n_35);
  L2_gameovercontrol_g3224 : AOI32D1BWP7T port map(A1 => L2_gameovercontrol_n_27, A2 => L2_gameovercontrol_n_3, A3 => L2_gameovercontrol_state(0), B1 => L2_gameovercontrol_n_21, B2 => L2_gameovercontrol_n_9, ZN => L2_gameovercontrol_n_34);
  L2_gameovercontrol_pixel_arr_buffer_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_30, Q => L2_gameovercontrol_pixel_arr_buffer(1));
  L2_gameovercontrol_pixel_arr_buffer_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_29, Q => L2_gameovercontrol_pixel_arr_buffer(2));
  L2_gameovercontrol_g3227 : MOAI22D0BWP7T port map(A1 => L2_gameovercontrol_n_24, A2 => L2_gameovercontrol_n_976_BAR, B1 => L2_gameovercontrol_n_27, B2 => L2_gameovercontrol_n_7, ZN => L2_gameovercontrol_n_32);
  L2_gameovercontrol_pixel_arr_buffer_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_28, Q => L2_gameovercontrol_pixel_arr_buffer(3));
  L2_gameovercontrol_g3230 : AO22D0BWP7T port map(A1 => L2_gameovercontrol_n_25, A2 => L2_gameovercontrol_pixel_arr_buffer(1), B1 => L2_gameovercontrol_n_26, B2 => L2_n_544, Z => L2_gameovercontrol_n_30);
  L2_gameovercontrol_g3231 : NR3D0BWP7T port map(A1 => L2_gameovercontrol_n_24, A2 => L2_gameovercontrol_state(0), A3 => L2_gameovercontrol_state(3), ZN => L2_gameovercontrol_n_31);
  L2_gameovercontrol_g3232 : AO22D0BWP7T port map(A1 => L2_gameovercontrol_n_25, A2 => L2_gameovercontrol_pixel_arr_buffer(2), B1 => L2_gameovercontrol_n_26, B2 => L2_n_540, Z => L2_gameovercontrol_n_29);
  L2_gameovercontrol_g3233 : AO22D0BWP7T port map(A1 => L2_gameovercontrol_n_25, A2 => L2_gameovercontrol_pixel_arr_buffer(3), B1 => L2_gameovercontrol_n_26, B2 => L2_n_541, Z => L2_gameovercontrol_n_28);
  L2_gameovercontrol_pixel_arr_buffer_reg_6 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_19, Q => L2_gameovercontrol_pixel_arr_buffer(6));
  L2_gameovercontrol_pixel_arr_buffer_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_23, Q => L2_gameovercontrol_pixel_arr_buffer(4));
  L2_gameovercontrol_pixel_arr_buffer_reg_5 : DFQD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_20, Q => L2_gameovercontrol_pixel_arr_buffer(5));
  L2_gameovercontrol_g3237 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_24, A2 => L2_gameovercontrol_n_10, ZN => L2_gameovercontrol_n_27);
  L2_gameovercontrol_g3238 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_18, A2 => reset, ZN => L2_gameovercontrol_n_26);
  L2_gameovercontrol_g3239 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_17, A2 => reset, ZN => L2_gameovercontrol_n_25);
  L2_gameovercontrol_g3241 : ND3D0BWP7T port map(A1 => L2_gameovercontrol_n_9, A2 => L2_gameovercontrol_n_164, A3 => L2_gameovercontrol_n_16, ZN => L2_gameovercontrol_n_24);
  L2_gameovercontrol_g3242 : AO22D0BWP7T port map(A1 => L2_n_542, A2 => L2_gameovercontrol_n_14, B1 => L2_gameovercontrol_pixel_arr_buffer(4), B2 => L2_gameovercontrol_n_15, Z => L2_gameovercontrol_n_23);
  L2_gameovercontrol_g3243 : OAI22D0BWP7T port map(A1 => L2_n_537, A2 => L2_gameovercontrol_n_16, B1 => L2_gameovercontrol_n_165, B2 => L2_gameovercontrol_n_164, ZN => L2_gameovercontrol_n_22);
  L2_gameovercontrol_g3244 : OAI22D0BWP7T port map(A1 => L2_gameovercontrol_n_4, A2 => L2_gameovercontrol_n_16, B1 => L2_gameovercontrol_n_5, B2 => L2_gameovercontrol_n_164, ZN => L2_gameovercontrol_n_21);
  L2_gameovercontrol_g3245 : AO22D0BWP7T port map(A1 => L2_n_543, A2 => L2_gameovercontrol_n_14, B1 => L2_gameovercontrol_pixel_arr_buffer(5), B2 => L2_gameovercontrol_n_15, Z => L2_gameovercontrol_n_20);
  L2_gameovercontrol_g3246 : AO22D0BWP7T port map(A1 => L2_n_545, A2 => L2_gameovercontrol_n_14, B1 => L2_gameovercontrol_pixel_arr_buffer(6), B2 => L2_gameovercontrol_n_15, Z => L2_gameovercontrol_n_19);
  L2_gameovercontrol_g3247 : CKND1BWP7T port map(I => L2_gameovercontrol_n_17, ZN => L2_gameovercontrol_n_18);
  L2_gameovercontrol_g3248 : OAI31D0BWP7T port map(A1 => L2_gameovercontrol_state(0), A2 => L2_gameovercontrol_n_3, A3 => L2_gameovercontrol_n_10, B => L2_gameovercontrol_n_13, ZN => L2_gameovercontrol_n_17);
  L2_gameovercontrol_g3249 : IND2D1BWP7T port map(A1 => L2_gameovercontrol_n_13, B1 => L2_gameovercontrol_state(0), ZN => L2_gameovercontrol_n_16);
  L2_gameovercontrol_g3250 : INR2D1BWP7T port map(A1 => L2_gameovercontrol_n_12, B1 => reset, ZN => L2_gameovercontrol_n_15);
  L2_gameovercontrol_g3251 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_n_12, A2 => reset, ZN => L2_gameovercontrol_n_14);
  L2_gameovercontrol_g3252 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_8, A2 => L2_gameovercontrol_n_3, ZN => L2_gameovercontrol_n_13);
  L2_gameovercontrol_g3253 : AOI21D0BWP7T port map(A1 => L2_gameovercontrol_n_162, A2 => L2_gameovercontrol_row, B => L2_gameovercontrol_n_2, ZN => L2_gameovercontrol_n_11);
  L2_gameovercontrol_g3254 : ND2D1BWP7T port map(A1 => L2_gameovercontrol_n_8, A2 => L2_gameovercontrol_n_7, ZN => L2_gameovercontrol_n_12);
  L2_gameovercontrol_g3255 : IND2D1BWP7T port map(A1 => L2_gameovercontrol_state(3), B1 => L2_gameovercontrol_state(2), ZN => L2_gameovercontrol_n_10);
  L2_gameovercontrol_g3256 : NR2D1BWP7T port map(A1 => L2_user_reset_new, A2 => reset, ZN => L2_gameovercontrol_n_9);
  L2_gameovercontrol_g3257 : INVD0BWP7T port map(I => L2_gameovercontrol_n_7, ZN => L2_gameovercontrol_n_6);
  L2_gameovercontrol_g3258 : NR2XD0BWP7T port map(A1 => L2_gameovercontrol_state(2), A2 => L2_gameovercontrol_state(3), ZN => L2_gameovercontrol_n_8);
  L2_gameovercontrol_g3259 : CKND2D1BWP7T port map(A1 => L2_gameovercontrol_state(0), A2 => L2_gameovercontrol_state(1), ZN => L2_gameovercontrol_n_7);
  L2_gameovercontrol_g3260 : INVD1BWP7T port map(I => L2_gameovercontrol_n_165, ZN => L2_gameovercontrol_n_5);
  L2_gameovercontrol_g3261 : INVD1BWP7T port map(I => L2_n_537, ZN => L2_gameovercontrol_n_4);
  L2_gameovercontrol_g3263 : INVD0BWP7T port map(I => L2_gameovercontrol_n_131, ZN => L2_gameovercontrol_n_2);
  L2_gameovercontrol_g2 : NR3D0BWP7T port map(A1 => L2_gameovercontrol_n_24, A2 => L2_gameovercontrol_n_163, A3 => L2_gameovercontrol_state(1), ZN => L2_gameovercontrol_n_166);
  L2_gameovercontrol_state_reg_3 : DFD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_35, Q => L2_gameovercontrol_state(3), QN => L2_gameovercontrol_n_45);
  L2_gameovercontrol_row_reg : DFXD1BWP7T port map(CP => clk, DA => L2_gameovercontrol_n_11, DB => L2_gameovercontrol_row, SA => L2_reset_county_go, Q => L2_gameovercontrol_row, QN => L2_gameovercontrol_n_40);
  L2_gameovercontrol_state_reg_1 : DFD1BWP7T port map(CP => clk, D => L2_gameovercontrol_n_36, Q => L2_gameovercontrol_state(1), QN => L2_gameovercontrol_n_3);
  L2_score_L2_in_c_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_score_L2_n_56, Q => L2_in_score_12bits(11));
  L2_score_L2_g1247 : OAI31D0BWP7T port map(A1 => L2_in_score_12bits(10), A2 => L2_score_L2_n_7, A3 => L2_score_L2_n_46, B => L2_score_L2_n_57, ZN => L2_score_L2_n_58);
  L2_score_L2_g1249 : OAI21D0BWP7T port map(A1 => L2_score_L2_n_50, A2 => L2_score_L2_n_36, B => L2_in_score_12bits(10), ZN => L2_score_L2_n_57);
  L2_score_L2_g1251 : OAI31D0BWP7T port map(A1 => L2_score_L2_n_7, A2 => L2_score_L2_n_4, A3 => L2_score_L2_n_46, B => L2_score_L2_n_53, ZN => L2_score_L2_n_56);
  L2_score_L2_g1252 : OAI221D0BWP7T port map(A1 => L2_score_L2_n_47, A2 => L2_score_L2_n_8, B1 => L2_in_score_12bits(8), B2 => L2_score_L2_n_41, C => L2_score_L2_n_51, ZN => L2_score_L2_n_55);
  L2_score_L2_in_b_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_score_L2_n_49, Q => L2_in_score_12bits(7));
  L2_score_L2_in_b_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_score_L2_n_48, Q => L2_in_score_12bits(5));
  L2_score_L2_g1255 : OAI21D0BWP7T port map(A1 => L2_score_L2_n_34, A2 => L2_in_score_12bits(6), B => L2_score_L2_n_52, ZN => L2_score_L2_n_54);
  L2_score_L2_g1256 : IOA21D1BWP7T port map(A1 => L2_score_L2_n_47, A2 => L2_score_L2_n_44, B => L2_in_score_12bits(11), ZN => L2_score_L2_n_53);
  L2_score_L2_g1257 : OAI21D0BWP7T port map(A1 => L2_score_L2_n_42, A2 => L2_score_L2_n_31, B => L2_in_score_12bits(6), ZN => L2_score_L2_n_52);
  L2_score_L2_g1258 : IND3D1BWP7T port map(A1 => L2_score_L2_n_44, B1 => L2_in_score_12bits(7), B2 => L2_score_L2_n_23, ZN => L2_score_L2_n_51);
  L2_score_L2_g1260 : MOAI22D0BWP7T port map(A1 => L2_score_L2_n_34, A2 => L2_score_L2_n_1, B1 => L2_score_L2_n_43, B2 => L2_in_score_12bits(7), ZN => L2_score_L2_n_49);
  L2_score_L2_g1261 : AO22D0BWP7T port map(A1 => L2_score_L2_n_42, A2 => L2_in_score_12bits(5), B1 => L2_score_L2_n_31, B2 => L2_score_L2_n_23, Z => L2_score_L2_n_48);
  L2_score_L2_g1262 : IOA21D1BWP7T port map(A1 => L2_score_L2_n_30, A2 => L2_score_L2_n_8, B => L2_score_L2_n_47, ZN => L2_score_L2_n_50);
  L2_score_L2_g1265 : INVD0BWP7T port map(I => L2_score_L2_n_45, ZN => L2_score_L2_n_46);
  L2_score_L2_g1266 : NR2XD0BWP7T port map(A1 => L2_score_L2_n_43, A2 => L2_score_L2_n_21, ZN => L2_score_L2_n_47);
  L2_score_L2_g1267 : NR2XD0BWP7T port map(A1 => L2_score_L2_n_41, A2 => L2_score_L2_n_8, ZN => L2_score_L2_n_45);
  L2_score_L2_g1269 : IND4D0BWP7T port map(A1 => L2_score_L2_n_24, B1 => L2_score_L2_n_7, B2 => L2_score_L2_n_4, B3 => L2_score_L2_n_8, ZN => L2_score_L2_n_44);
  L2_score_L2_g1270 : AOI21D0BWP7T port map(A1 => L2_score_L2_n_27, A2 => L2_score_L2_n_19, B => L2_score_reset_or, ZN => L2_score_L2_n_43);
  L2_score_L2_g1271 : AO21D0BWP7T port map(A1 => L2_score_L2_n_21, A2 => L2_score_L2_n_0, B => L2_score_L2_n_37, Z => L2_score_L2_n_42);
  L2_score_L2_in_a_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_score_L2_n_32, Q => L2_in_score_12bits(1));
  L2_score_L2_g1273 : OAI22D0BWP7T port map(A1 => L2_score_L2_n_28, A2 => L2_score_L2_n_9, B1 => L2_score_L2_n_29, B2 => L2_score_reset_or, ZN => L2_score_L2_n_40);
  L2_score_L2_g1274 : OAI31D0BWP7T port map(A1 => L2_score_L2_n_5, A2 => L2_score_reset_or, A3 => score_pulse_int, B => L2_score_L2_n_35, ZN => L2_score_L2_n_39);
  L2_score_L2_g1275 : MOAI22D0BWP7T port map(A1 => L2_score_L2_n_28, A2 => L2_in_score_12bits(2), B1 => L2_score_L2_n_26, B2 => L2_in_score_12bits(2), ZN => L2_score_L2_n_38);
  L2_score_L2_g1276 : ND3D0BWP7T port map(A1 => L2_score_L2_n_23, A2 => L2_score_L2_n_30, A3 => L2_in_score_12bits(7), ZN => L2_score_L2_n_41);
  L2_score_L2_g1277 : AN2D0BWP7T port map(A1 => L2_score_L2_n_30, A2 => L2_score_L2_n_7, Z => L2_score_L2_n_36);
  L2_score_L2_g1278 : OAI211D1BWP7T port map(A1 => L2_score_L2_n_10, A2 => L2_score_L2_n_16, B => score_pulse_int, C => L2_score_L2_n_5, ZN => L2_score_L2_n_35);
  L2_score_L2_g1279 : NR2D1BWP7T port map(A1 => L2_score_L2_n_27, A2 => L2_score_reset_or, ZN => L2_score_L2_n_37);
  L2_score_L2_g1280 : AOI21D0BWP7T port map(A1 => L2_score_L2_n_20, A2 => L2_score_L2_n_24, B => L2_score_L2_n_17, ZN => L2_score_L2_n_33);
  L2_score_L2_g1281 : AO22D0BWP7T port map(A1 => L2_score_L2_n_18, A2 => L2_score_L2_n_11, B1 => L2_in_score_12bits(1), B2 => L2_score_L2_n_25, Z => L2_score_L2_n_32);
  L2_score_L2_g1282 : ND3D0BWP7T port map(A1 => L2_score_L2_n_23, A2 => L2_score_L2_n_21, A3 => L2_in_score_12bits(5), ZN => L2_score_L2_n_34);
  L2_score_L2_g1283 : ND2D1BWP7T port map(A1 => L2_score_L2_n_22, A2 => L2_in_score_12bits(3), ZN => L2_score_L2_n_29);
  L2_score_L2_g1284 : NR2D1BWP7T port map(A1 => L2_score_L2_n_20, A2 => L2_in_score_12bits(5), ZN => L2_score_L2_n_31);
  L2_score_L2_g1285 : NR2XD0BWP7T port map(A1 => L2_score_L2_n_24, A2 => L2_in_score_12bits(11), ZN => L2_score_L2_n_30);
  L2_score_L2_g1286 : AO21D0BWP7T port map(A1 => L2_score_L2_n_11, A2 => L2_score_L2_n_6, B => L2_score_L2_n_25, Z => L2_score_L2_n_26);
  L2_score_L2_g1287 : IND3D1BWP7T port map(A1 => L2_score_reset_or, B1 => L2_in_score_12bits(1), B2 => L2_score_L2_n_18, ZN => L2_score_L2_n_28);
  L2_score_L2_g1288 : INR2XD0BWP7T port map(A1 => L2_in_score_12bits(3), B1 => L2_score_L2_n_22, ZN => L2_score_L2_n_27);
  L2_score_L2_g1289 : AOI21D0BWP7T port map(A1 => score_pulse_int, A2 => L2_score_L2_n_13, B => L2_score_reset_or, ZN => L2_score_L2_n_25);
  L2_score_L2_g1290 : ND2D1BWP7T port map(A1 => L2_score_L2_n_16, A2 => L2_score_L2_n_12, ZN => L2_score_L2_n_24);
  L2_score_L2_g1291 : NR2XD0BWP7T port map(A1 => L2_score_L2_n_17, A2 => L2_score_L2_n_0, ZN => L2_score_L2_n_23);
  L2_score_L2_g1292 : INVD0BWP7T port map(I => L2_score_L2_n_21, ZN => L2_score_L2_n_20);
  L2_score_L2_g1293 : ND3D0BWP7T port map(A1 => L2_score_L2_n_14, A2 => L2_score_L2_n_12, A3 => L2_score_L2_n_0, ZN => L2_score_L2_n_19);
  L2_score_L2_g1294 : IOA21D1BWP7T port map(A1 => L2_score_L2_n_14, A2 => L2_score_L2_n_5, B => score_pulse_int, ZN => L2_score_L2_n_22);
  L2_score_L2_g1295 : INR2D1BWP7T port map(A1 => L2_score_L2_n_16, B1 => L2_in_score_12bits(7), ZN => L2_score_L2_n_21);
  L2_score_L2_g1296 : NR2XD0BWP7T port map(A1 => L2_score_L2_n_15, A2 => L2_in_score_12bits(3), ZN => L2_score_L2_n_18);
  L2_score_L2_g1297 : OR2D1BWP7T port map(A1 => L2_score_L2_n_15, A2 => L2_score_L2_n_6, Z => L2_score_L2_n_17);
  L2_score_L2_g1298 : CKAN2D1BWP7T port map(A1 => L2_score_L2_n_11, A2 => L2_score_L2_n_9, Z => L2_score_L2_n_16);
  L2_score_L2_g1299 : ND2D1BWP7T port map(A1 => L2_score_L2_n_5, A2 => L2_score_L2_n_6, ZN => L2_score_L2_n_13);
  L2_score_L2_g1300 : ND2D1BWP7T port map(A1 => score_pulse_int, A2 => L2_in_score_12bits(0), ZN => L2_score_L2_n_15);
  L2_score_L2_g1301 : NR2XD0BWP7T port map(A1 => L2_in_score_12bits(1), A2 => L2_in_score_12bits(2), ZN => L2_score_L2_n_14);
  L2_score_L2_g1302 : NR2XD0BWP7T port map(A1 => L2_score_reset_or, A2 => L2_in_score_12bits(3), ZN => L2_score_L2_n_10);
  L2_score_L2_g1303 : NR2XD0BWP7T port map(A1 => L2_in_score_12bits(5), A2 => L2_in_score_12bits(6), ZN => L2_score_L2_n_12);
  L2_score_L2_g1304 : NR2XD0BWP7T port map(A1 => L2_score_reset_or, A2 => L2_in_score_12bits(1), ZN => L2_score_L2_n_11);
  L2_score_L2_in_c_reg_2 : DFD1BWP7T port map(CP => clk, D => L2_score_L2_n_58, Q => L2_in_score_12bits(10), QN => L2_score_L2_n_4);
  L2_score_L2_in_a_reg_2 : DFD1BWP7T port map(CP => clk, D => L2_score_L2_n_38, Q => L2_in_score_12bits(2), QN => L2_score_L2_n_9);
  L2_score_L2_in_c_reg_0 : DFD1BWP7T port map(CP => clk, D => L2_score_L2_n_55, Q => L2_in_score_12bits(8), QN => L2_score_L2_n_8);
  L2_score_L2_in_c_reg_1 : DFXD1BWP7T port map(CP => clk, DA => L2_score_L2_n_50, DB => L2_score_L2_n_45, SA => L2_in_score_12bits(9), Q => L2_in_score_12bits(9), QN => L2_score_L2_n_7);
  L2_score_L2_in_a_reg_3 : DFD1BWP7T port map(CP => clk, D => L2_score_L2_n_40, Q => L2_in_score_12bits(3), QN => L2_score_L2_n_6);
  L2_score_L2_in_b_reg_2 : DFD1BWP7T port map(CP => clk, D => L2_score_L2_n_54, Q => L2_in_score_12bits(6), QN => L2_score_L2_n_1);
  L2_score_L2_in_a_reg_0 : DFD1BWP7T port map(CP => clk, D => L2_score_L2_n_39, Q => L2_in_score_12bits(0), QN => L2_score_L2_n_5);
  L2_score_L2_in_b_reg_0 : DFXD1BWP7T port map(CP => clk, DA => L2_score_L2_n_37, DB => L2_score_L2_n_33, SA => L2_in_score_12bits(4), Q => L2_in_score_12bits(4), QN => L2_score_L2_n_0);
  L2_score_L3_score_type_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_81, Q => L2_score_score_sprite_type(0));
  L2_score_L3_score_type_reg_1 : DFQD0BWP7T port map(CP => clk, D => L2_score_L3_n_80, Q => L2_score_score_sprite_type(1));
  L2_score_L3_score_type_reg_2 : DFQD0BWP7T port map(CP => clk, D => L2_score_L3_n_79, Q => L2_score_score_sprite_type(2));
  L2_score_L3_score_type_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_78, Q => L2_score_score_sprite_type(3));
  L2_score_L3_g2368 : AO221D0BWP7T port map(A1 => L2_score_L3_n_66, A2 => L2_in_score_12bits(4), B1 => L2_score_L3_n_68, B2 => L2_in_score_12bits(0), C => L2_score_L3_n_77, Z => L2_score_L3_n_81);
  L2_score_L3_g2369 : ND2D1BWP7T port map(A1 => L2_score_L3_n_76, A2 => L2_score_L3_n_73, ZN => L2_score_L3_n_80);
  L2_score_L3_g2370 : AO221D0BWP7T port map(A1 => L2_score_L3_n_66, A2 => L2_in_score_12bits(6), B1 => L2_score_L3_n_69, B2 => L2_in_score_12bits(10), C => L2_score_L3_n_74, Z => L2_score_L3_n_79);
  L2_score_L3_g2371 : AO221D0BWP7T port map(A1 => L2_score_L3_n_66, A2 => L2_in_score_12bits(7), B1 => L2_score_L3_n_69, B2 => L2_in_score_12bits(11), C => L2_score_L3_n_75, Z => L2_score_L3_n_78);
  L2_score_L3_g2372 : OAI21D0BWP7T port map(A1 => L2_score_L3_n_72, A2 => L2_score_L3_n_41, B => L2_score_L3_n_48, ZN => L2_reset_county_score);
  L2_score_L3_g2373 : OAI31D0BWP7T port map(A1 => L2_current_block_horizontal(0), A2 => L2_score_L3_n_51, A3 => L2_score_L3_n_67, B => L2_score_L3_n_71, ZN => L2_score_L3_n_77);
  L2_score_L3_g2374 : INR2XD0BWP7T port map(A1 => L2_score_L3_n_41, B1 => L2_score_L3_n_72, ZN => L2_en_county_score);
  L2_score_L3_g2375 : ND2D1BWP7T port map(A1 => L2_score_L3_n_72, A2 => L2_score_L3_n_48, ZN => L2_reset_dual_pixel_y_score);
  L2_score_L3_g2376 : IND3D1BWP7T port map(A1 => L2_score_L3_n_93, B1 => L2_score_L3_n_83, B2 => L2_score_L3_n_65, ZN => L2_rgb_score(0));
  L2_score_L3_g2377 : AOI22D0BWP7T port map(A1 => L2_score_L3_n_66, A2 => L2_in_score_12bits(5), B1 => L2_score_L3_n_69, B2 => L2_in_score_12bits(9), ZN => L2_score_L3_n_76);
  L2_score_L3_g2378 : MOAI22D0BWP7T port map(A1 => L2_score_L3_n_67, A2 => L2_score_L3_n_52, B1 => L2_score_L3_n_68, B2 => L2_in_score_12bits(3), ZN => L2_score_L3_n_75);
  L2_score_L3_g2379 : MOAI22D0BWP7T port map(A1 => L2_score_L3_n_67, A2 => L2_score_L3_n_53, B1 => L2_score_L3_n_68, B2 => L2_in_score_12bits(2), ZN => L2_score_L3_n_74);
  L2_score_L3_g2380 : MAOI22D0BWP7T port map(A1 => L2_score_L3_n_68, A2 => L2_in_score_12bits(1), B1 => L2_score_L3_n_67, B2 => L2_score_L3_n_57, ZN => L2_score_L3_n_73);
  L2_score_L3_g2381 : IND2D1BWP7T port map(A1 => L2_score_L3_n_70, B1 => L2_score_L3_n_48, ZN => L2_reset_current_block_horizontal_score);
  L2_score_L3_g2382 : INR2D1BWP7T port map(A1 => L2_score_L3_n_70, B1 => L2_dual_pixel_y, ZN => L2_en_dual_pixel_y_score);
  L2_score_L3_g2383 : ND2D1BWP7T port map(A1 => L2_score_L3_n_69, A2 => L2_in_score_12bits(8), ZN => L2_score_L3_n_71);
  L2_score_L3_g2384 : ND2D1BWP7T port map(A1 => L2_score_L3_n_70, A2 => L2_dual_pixel_y, ZN => L2_score_L3_n_72);
  L2_score_L3_g2385 : INR2XD0BWP7T port map(A1 => L2_score_L3_n_135, B1 => L2_score_L3_n_83, ZN => L2_en_current_block_horizontal_score);
  L2_score_L3_g2386 : NR2D1BWP7T port map(A1 => L2_score_L3_n_135, A2 => L2_score_L3_n_83, ZN => L2_score_L3_n_70);
  L2_score_L3_g2387 : AN2D1BWP7T port map(A1 => L2_score_L3_n_30, A2 => L2_score_L3_n_45, Z => L2_score_L3_n_69);
  L2_score_L3_g2388 : INR2D1BWP7T port map(A1 => L2_score_L3_n_30, B1 => L2_score_L3_n_45, ZN => L2_score_L3_n_68);
  L2_score_L3_g2389 : ND3D0BWP7T port map(A1 => L2_score_L3_n_61, A2 => L2_score_L3_n_60, A3 => L2_score_L3_n_56, ZN => L2_rgb_score(2));
  L2_score_L3_g2390 : NR3D0BWP7T port map(A1 => L2_score_L3_n_55, A2 => L2_score_L3_n_59, A3 => L2_score_L3_n_62, ZN => L2_score_L3_n_65);
  L2_score_L3_g2391 : ND2D1BWP7T port map(A1 => L2_score_L3_n_63, A2 => L2_score_L3_n_45, ZN => L2_score_L3_n_67);
  L2_score_L3_g2392 : NR2D1BWP7T port map(A1 => L2_score_L3_n_64, A2 => L2_score_L3_n_45, ZN => L2_score_L3_n_66);
  L2_score_L3_g2393 : OAI21D0BWP7T port map(A1 => L2_score_L3_n_54, A2 => L2_current_block_horizontal(3), B => L2_current_block_horizontal(4), ZN => L2_score_L3_n_135);
  L2_score_L3_g2394 : INVD0BWP7T port map(I => L2_score_L3_n_63, ZN => L2_score_L3_n_64);
  L2_score_L3_g2396 : NR2D1BWP7T port map(A1 => L2_score_reset_or, A2 => L2_score_L3_n_58, ZN => L2_score_L3_n_63);
  L2_score_L3_g2397 : OAI33D1BWP7T port map(A1 => L2_score_L3_pixel_arr_buffer(2), A2 => L2_score_L3_state(1), A3 => L2_score_L3_n_44, B1 => L2_score_L3_pixel_arr_buffer(3), B2 => L2_score_L3_state(1), B3 => L2_score_L3_n_29, ZN => L2_score_L3_n_62);
  L2_score_L3_g2398 : AOI22D0BWP7T port map(A1 => L2_score_L3_n_90, A2 => L2_score_L3_pixel_arr_buffer(2), B1 => L2_score_L3_n_89, B2 => L2_score_L3_pixel_arr_buffer(3), ZN => L2_score_L3_n_61);
  L2_score_L3_g2399 : AOI22D0BWP7T port map(A1 => L2_score_L3_n_2, A2 => L2_score_L3_pixel_arr_buffer(4), B1 => L2_score_L3_n_88, B2 => L2_score_L3_pixel_arr_buffer(5), ZN => L2_score_L3_n_60);
  L2_score_L3_g2400 : OAI22D0BWP7T port map(A1 => L2_score_L3_n_46, A2 => L2_score_L3_pixel_arr_buffer(4), B1 => L2_score_L3_n_50, B2 => L2_score_L3_pixel_arr_buffer(5), ZN => L2_score_L3_n_59);
  L2_score_L3_g2402 : MAOI22D0BWP7T port map(A1 => L2_score_L3_n_42, A2 => L2_score_L3_n_35, B1 => L2_score_L3_n_40, B2 => L2_score_L3_n_39, ZN => L2_score_L3_n_57);
  L2_score_L3_g2403 : AOI22D0BWP7T port map(A1 => L2_score_L3_n_87, A2 => L2_score_L3_pixel_arr_buffer(6), B1 => L2_score_L3_n_91, B2 => L2_score_L3_pixel_arr_buffer(1), ZN => L2_score_L3_n_56);
  L2_score_L3_g2404 : OAI22D0BWP7T port map(A1 => L2_score_L3_n_47, A2 => L2_score_L3_pixel_arr_buffer(6), B1 => L2_score_L3_n_49, B2 => L2_score_L3_pixel_arr_buffer(1), ZN => L2_score_L3_n_55);
  L2_score_L3_g2405 : OAI22D0BWP7T port map(A1 => L2_score_L3_n_45, A2 => L2_score_L3_n_31, B1 => L2_score_L3_n_43, B2 => L2_score_L3_n_33, ZN => L2_score_L3_n_58);
  L2_score_L3_g2406 : INR2D1BWP7T port map(A1 => L2_current_block_horizontal(2), B1 => L2_score_L3_n_33, ZN => L2_score_L3_n_54);
  L2_score_L3_g2407 : INR2XD0BWP7T port map(A1 => L2_score_L3_n_35, B1 => L2_score_L3_n_40, ZN => L2_score_L3_n_53);
  L2_score_L3_g2408 : NR2XD0BWP7T port map(A1 => L2_score_L3_n_40, A2 => L2_score_L3_n_33, ZN => L2_score_L3_n_52);
  L2_score_L3_g2409 : OA21D0BWP7T port map(A1 => L2_score_L3_n_40, A2 => L2_score_L3_n_32, B => L2_score_L3_n_43, Z => L2_score_L3_n_51);
  L2_score_L3_g2410 : INVD0BWP7T port map(I => L2_score_L3_n_88, ZN => L2_score_L3_n_50);
  L2_score_L3_g2411 : INVD1BWP7T port map(I => L2_score_L3_n_49, ZN => L2_score_L3_n_91);
  L2_score_L3_g2412 : NR2D1BWP7T port map(A1 => L2_score_L3_n_44, A2 => L2_score_L3_state(1), ZN => L2_score_L3_n_90);
  L2_score_L3_g2413 : INR2D1BWP7T port map(A1 => L2_score_L3_state(1), B1 => L2_score_L3_n_29, ZN => L2_score_L3_n_88);
  L2_score_L3_g2414 : NR2D1BWP7T port map(A1 => L2_score_L3_n_29, A2 => L2_score_L3_state(1), ZN => L2_score_L3_n_89);
  L2_score_L3_g2415 : ND2D1BWP7T port map(A1 => L2_score_L3_n_94, A2 => L2_score_L3_state(1), ZN => L2_score_L3_n_49);
  L2_score_L3_g2416 : INR2XD0BWP7T port map(A1 => L2_score_L3_n_84, B1 => L2_score_L3_n_95, ZN => L2_score_L3_n_48);
  L2_score_L3_g2417 : INVD1BWP7T port map(I => L2_score_L3_n_47, ZN => L2_score_L3_n_87);
  L2_score_L3_g2418 : INVD0BWP7T port map(I => L2_score_L3_n_2, ZN => L2_score_L3_n_46);
  L2_score_L3_g2420 : IND3D0BWP7T port map(A1 => L2_score_L3_state(0), B1 => L2_score_L3_state(3), B2 => L2_score_L3_n_36, ZN => L2_score_L3_n_47);
  L2_score_L3_g2421 : INR2D1BWP7T port map(A1 => L2_score_L3_state(1), B1 => L2_score_L3_n_44, ZN => L2_score_L3_n_2);
  L2_score_L3_g2422 : ND3D0BWP7T port map(A1 => L2_score_L3_n_36, A2 => L2_score_L3_state(3), A3 => L2_score_L3_state(0), ZN => L2_score_L3_n_83);
  L2_score_L3_g2423 : ND3D0BWP7T port map(A1 => L2_score_L3_n_38, A2 => L2_score_L3_n_32, A3 => L2_current_block_horizontal(2), ZN => L2_score_L3_n_45);
  L2_score_L3_g2424 : INVD0BWP7T port map(I => L2_score_L3_n_43, ZN => L2_score_L3_n_42);
  L2_score_L3_g2425 : IND2D1BWP7T port map(A1 => L2_score_L3_n_37, B1 => L2_score_L3_state(2), ZN => L2_score_L3_n_44);
  L2_score_L3_g2426 : NR2XD0BWP7T port map(A1 => L2_score_L3_n_34, A2 => L2_score_L3_state(2), ZN => L2_score_L3_n_94);
  L2_score_L3_g2428 : IND2D1BWP7T port map(A1 => L2_current_block_horizontal(2), B1 => L2_score_L3_n_38, ZN => L2_score_L3_n_43);
  L2_score_L3_g2429 : AOI22D0BWP7T port map(A1 => L2_score_L3_n_31, A2 => L2_current_block_horizontal(1), B1 => L2_score_L3_n_32, B2 => L2_current_block_horizontal(0), ZN => L2_score_L3_n_39);
  L2_score_L3_g2430 : IND2D1BWP7T port map(A1 => L2_score_L3_n_36, B1 => L2_score_L3_state(3), ZN => L2_score_L3_n_84);
  L2_score_L3_g2431 : INR2D1BWP7T port map(A1 => L2_score_L3_n_36, B1 => L2_score_L3_n_37, ZN => L2_score_L3_n_95);
  L2_score_L3_g2432 : ND3D0BWP7T port map(A1 => L2_county(2), A2 => L2_in_go_y_pos(1), A3 => L2_county(0), ZN => L2_score_L3_n_41);
  L2_score_L3_g2433 : IND3D1BWP7T port map(A1 => L2_current_block_horizontal(4), B1 => L2_current_block_horizontal(3), B2 => L2_current_block_horizontal(2), ZN => L2_score_L3_n_40);
  L2_score_L3_g2434 : INR2XD0BWP7T port map(A1 => L2_current_block_horizontal(4), B1 => L2_current_block_horizontal(3), ZN => L2_score_L3_n_38);
  L2_score_L3_g2435 : OR2D1BWP7T port map(A1 => L2_score_L3_state(3), A2 => L2_score_L3_state(0), Z => L2_score_L3_n_37);
  L2_score_L3_g2436 : NR2XD0BWP7T port map(A1 => L2_score_L3_state(1), A2 => L2_score_L3_state(2), ZN => L2_score_L3_n_36);
  L2_score_L3_g2438 : CKND2D1BWP7T port map(A1 => L2_score_L3_n_32, A2 => L2_score_L3_n_31, ZN => L2_score_L3_n_35);
  L2_score_L3_g2439 : IND2D1BWP7T port map(A1 => L2_score_L3_state(3), B1 => L2_score_L3_state(0), ZN => L2_score_L3_n_34);
  L2_score_L3_g2440 : CKND2D1BWP7T port map(A1 => L2_current_block_horizontal(1), A2 => L2_current_block_horizontal(0), ZN => L2_score_L3_n_33);
  L2_score_L3_g2441 : INVD1BWP7T port map(I => L2_current_block_horizontal(1), ZN => L2_score_L3_n_32);
  L2_score_L3_g2442 : INVD0BWP7T port map(I => L2_current_block_horizontal(0), ZN => L2_score_L3_n_31);
  L2_score_L3_g2 : INR2D1BWP7T port map(A1 => L2_score_L3_n_58, B1 => L2_score_reset_or, ZN => L2_score_L3_n_30);
  L2_score_L3_g2444 : IND2D1BWP7T port map(A1 => L2_score_L3_n_34, B1 => L2_score_L3_state(2), ZN => L2_score_L3_n_29);
  L2_score_L3_g2445 : INR3D0BWP7T port map(A1 => L2_score_L3_state(1), B1 => L2_score_L3_n_37, B2 => L2_score_L3_state(2), ZN => L2_score_L3_n_93);
  L2_score_L3_pixel_arr_buffer_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_27, Q => L2_score_L3_pixel_arr_buffer(1));
  L2_score_L3_pixel_arr_buffer_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_28, Q => L2_score_L3_pixel_arr_buffer(2));
  L2_score_L3_pixel_arr_buffer_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_26, Q => L2_score_L3_pixel_arr_buffer(3));
  L2_score_L3_pixel_arr_buffer_reg_5 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_22, Q => L2_score_L3_pixel_arr_buffer(5));
  L2_score_L3_pixel_arr_buffer_reg_6 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_24, Q => L2_score_L3_pixel_arr_buffer(6));
  L2_score_L3_pixel_arr_buffer_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_23, Q => L2_score_L3_pixel_arr_buffer(4));
  L2_score_L3_g1660 : AO22D0BWP7T port map(A1 => L2_score_L3_n_20, A2 => L2_score_L3_pixel_arr_buffer(2), B1 => L2_score_L3_n_15, B2 => L2_n_546, Z => L2_score_L3_n_28);
  L2_score_L3_g1661 : AO22D0BWP7T port map(A1 => L2_score_L3_n_20, A2 => L2_score_L3_pixel_arr_buffer(1), B1 => L2_score_L3_n_15, B2 => L2_n_550, Z => L2_score_L3_n_27);
  L2_score_L3_g1662 : AO22D0BWP7T port map(A1 => L2_score_L3_n_20, A2 => L2_score_L3_pixel_arr_buffer(3), B1 => L2_score_L3_n_15, B2 => L2_n_547, Z => L2_score_L3_n_26);
  L2_score_L3_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_25, Q => L2_score_L3_state(1));
  L2_score_L3_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_19, Q => L2_score_L3_state(0));
  L2_score_L3_state_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_score_L3_n_21, Q => L2_score_L3_state(2));
  L2_score_L3_g1666 : AO221D0BWP7T port map(A1 => L2_score_L3_n_8, A2 => L2_score_L3_n_5, B1 => L2_score_L3_n_9, B2 => L2_score_L3_n_93, C => L2_score_L3_n_16, Z => L2_score_L3_n_25);
  L2_score_L3_g1667 : AO22D0BWP7T port map(A1 => L2_score_L3_n_17, A2 => L2_score_L3_pixel_arr_buffer(6), B1 => L2_score_L3_n_18, B2 => L2_n_551, Z => L2_score_L3_n_24);
  L2_score_L3_g1668 : AO22D0BWP7T port map(A1 => L2_score_L3_n_17, A2 => L2_score_L3_pixel_arr_buffer(4), B1 => L2_score_L3_n_18, B2 => L2_n_548, Z => L2_score_L3_n_23);
  L2_score_L3_g1669 : AO22D0BWP7T port map(A1 => L2_score_L3_n_17, A2 => L2_score_L3_pixel_arr_buffer(5), B1 => L2_n_549, B2 => L2_score_L3_n_18, Z => L2_score_L3_n_22);
  L2_score_L3_state_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_score_L3_n_1, D => L2_score_L3_n_9, Q => L2_score_L3_state(3));
  L2_score_L3_g1671 : IND2D1BWP7T port map(A1 => L2_score_L3_n_16, B1 => L2_score_L3_n_14, ZN => L2_score_L3_n_21);
  L2_score_L3_g1672 : AO22D0BWP7T port map(A1 => L2_score_L3_n_9, A2 => L2_score_L3_n_10, B1 => L2_score_L3_n_5, B2 => L2_score_L3_n_7, Z => L2_score_L3_n_19);
  L2_score_L3_g1673 : NR3D0BWP7T port map(A1 => L2_score_reset_or, A2 => L2_score_L3_n_6, A3 => L2_score_L3_n_2, ZN => L2_score_L3_n_20);
  L2_score_L3_g1674 : NR2D1BWP7T port map(A1 => L2_score_reset_or, A2 => L2_score_L3_n_12, ZN => L2_score_L3_n_18);
  L2_score_L3_g1675 : NR2D1BWP7T port map(A1 => L2_score_reset_or, A2 => L2_score_L3_n_13, ZN => L2_score_L3_n_17);
  L2_score_L3_g1676 : OAI21D0BWP7T port map(A1 => L2_score_L3_n_91, A2 => L2_score_L3_n_90, B => L2_score_L3_n_9, ZN => L2_score_L3_n_14);
  L2_score_L3_g1677 : OA21D0BWP7T port map(A1 => L2_score_L3_n_89, A2 => L2_score_L3_n_2, B => L2_score_L3_n_9, Z => L2_score_L3_n_16);
  L2_score_L3_g1678 : IAO21D0BWP7T port map(A1 => L2_score_L3_n_2, A2 => L2_score_L3_n_6, B => L2_score_reset_or, ZN => L2_score_L3_n_15);
  L2_score_L3_g1679 : INVD0BWP7T port map(I => L2_score_L3_n_12, ZN => L2_score_L3_n_13);
  L2_score_L3_g1681 : INR4D0BWP7T port map(A1 => L2_score_L3_n_84, B1 => L2_score_L3_n_89, B2 => L2_score_L3_n_91, B3 => L2_score_L3_n_88, ZN => L2_score_L3_n_10);
  L2_score_L3_g1682 : NR2XD0BWP7T port map(A1 => L2_score_L3_n_6, A2 => L2_score_L3_n_93, ZN => L2_score_L3_n_12);
  L2_score_L3_g1683 : MOAI22D0BWP7T port map(A1 => L2_score_L3_n_0, A2 => L2_score_L3_n_83, B1 => L2_n_535, B2 => L2_score_L3_n_3, ZN => L2_score_L3_n_8);
  L2_score_L3_g1684 : OAI22D0BWP7T port map(A1 => L2_n_535, A2 => L2_score_L3_n_4, B1 => L2_score_L3_n_135, B2 => L2_score_L3_n_83, ZN => L2_score_L3_n_7);
  L2_score_L3_g1685 : AN3D1BWP7T port map(A1 => L2_score_L3_n_5, A2 => L2_score_L3_n_4, A3 => L2_score_L3_n_83, Z => L2_score_L3_n_9);
  L2_score_L3_g1686 : IND2D1BWP7T port map(A1 => L2_score_L3_n_95, B1 => L2_score_L3_n_4, ZN => L2_score_L3_n_6);
  L2_score_L3_g1687 : INVD0BWP7T port map(I => L2_score_L3_n_4, ZN => L2_score_L3_n_3);
  L2_score_L3_g1688 : NR2D1BWP7T port map(A1 => L2_user_reset_new, A2 => L2_score_reset_or, ZN => L2_score_L3_n_5);
  L2_score_L3_g1689 : IND2D1BWP7T port map(A1 => L2_score_L3_state(1), B1 => L2_score_L3_n_94, ZN => L2_score_L3_n_4);
  L2_score_L3_g1690 : OR2D1BWP7T port map(A1 => L2_score_L3_n_88, A2 => L2_score_L3_n_87, Z => L2_score_L3_n_1);
  L2_score_L3_g1692 : CKND1BWP7T port map(I => L2_score_L3_n_135, ZN => L2_score_L3_n_0);
  L2_shift_L11_g12367 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_276, A2 => L2_county(0), B => L2_shift_L11_n_285, ZN => L2_shift_y_pos_out_shift_pacman(0));
  L2_shift_L11_g12368 : OR4D1BWP7T port map(A1 => L2_shift_L11_n_256, A2 => L2_shift_L11_n_272, A3 => L2_shift_L11_n_275, A4 => L2_shift_L11_n_283, Z => L2_shift_y_pos_out_shift_pacman(2));
  L2_shift_L11_g12369 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_173, A2 => L2_shift_L11_n_144, B => L2_shift_L11_n_284, C => L2_shift_L11_n_274, ZN => L2_shift_y_pos_out_shift_pacman(1));
  L2_shift_L11_g12370 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_282, A2 => L2_shift_L11_n_269, B => L2_county(0), ZN => L2_shift_L11_n_285);
  L2_shift_L11_g12371 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_282, A2 => L2_in_go_y_pos(1), B1 => L2_shift_L11_n_270, B2 => L2_shift_L11_n_173, ZN => L2_shift_L11_n_284);
  L2_shift_L11_g12372 : MOAI22D0BWP7T port map(A1 => L2_shift_L11_n_267, A2 => L2_shift_L11_n_175, B1 => L2_shift_L11_n_281, B2 => L2_county(2), ZN => L2_shift_L11_n_283);
  L2_shift_L11_g12373 : OR2D1BWP7T port map(A1 => L2_shift_L11_n_281, A2 => L2_shift_L11_n_290, Z => L2_shift_L11_n_282);
  L2_shift_L11_g12374 : IND2D1BWP7T port map(A1 => L2_shift_cell_state_out_shift_pacman(4), B1 => L2_shift_L11_n_280, ZN => L2_n_531);
  L2_shift_L11_g12375 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_278, A2 => L2_shift_L11_n_289, A3 => L2_shift_L11_n_293, A4 => L2_shift_L11_n_290, ZN => L2_shift_L11_n_281);
  L2_shift_L11_g12376 : AOI211XD0BWP7T port map(A1 => L2_shift_L11_n_260, A2 => L2_shift_L11_n_307, B => cell_type_int(0), C => L2_shift_L11_n_279, ZN => L2_shift_L11_n_280);
  L2_shift_L11_g12377 : CKAN2D1BWP7T port map(A1 => cell_type_int(1), A2 => L2_shift_L11_n_277, Z => L2_shift_cell_state_out_shift_pacman(1));
  L2_shift_L11_g12378 : AN2D1BWP7T port map(A1 => cell_type_int(2), A2 => L2_shift_L11_n_277, Z => L2_shift_cell_state_out_shift_pacman(2));
  L2_shift_L11_g12379 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_271, A2 => L2_shift_L11_n_260, A3 => L2_shift_L11_n_230, A4 => L2_shift_L11_n_214, ZN => L2_shift_L11_n_279);
  L2_shift_L11_g12380 : OR4XD1BWP7T port map(A1 => L2_shift_L11_n_287, A2 => L2_shift_L11_n_264, A3 => L2_shift_L11_n_269, A4 => L2_shift_L11_n_270, Z => L2_shift_L11_n_278);
  L2_shift_L11_g12381 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_271, B1 => L2_shift_L11_n_273, ZN => L2_shift_L11_n_277);
  L2_shift_L11_g12382 : INR2XD0BWP7T port map(A1 => L2_shift_L11_n_144, B1 => L2_shift_L11_n_270, ZN => L2_shift_L11_n_276);
  L2_shift_L11_g12383 : AO222D0BWP7T port map(A1 => L2_shift_L11_n_266, A2 => L2_shift_L11_n_203, B1 => L2_shift_L11_n_263, B2 => L2_shift_L11_n_175, C1 => L2_shift_L11_n_264, C2 => L2_shift_L11_n_212, Z => L2_shift_L11_n_275);
  L2_shift_L11_g12384 : AO21D0BWP7T port map(A1 => L2_shift_L11_n_267, A2 => L2_shift_L11_n_262, B => L2_in_go_y_pos(1), Z => L2_shift_L11_n_274);
  L2_shift_L11_g12386 : AOI222D0BWP7T port map(A1 => L2_shift_L11_n_260, A2 => L2_shift_L11_n_227, B1 => L2_shift_L11_n_296, B2 => L2_shift_L11_n_230, C1 => L2_shift_L11_n_298, C2 => L2_shift_L11_n_214, ZN => L2_shift_L11_n_273);
  L2_shift_L11_g12387 : OAI22D0BWP7T port map(A1 => L2_shift_L11_n_268, A2 => L2_shift_L11_n_212, B1 => L2_shift_L11_n_265, B2 => L2_shift_L11_n_203, ZN => L2_shift_L11_n_272);
  L2_shift_L11_g12388 : AO221D0BWP7T port map(A1 => L2_shift_L11_n_297, A2 => L2_shift_L11_n_210, B1 => L2_shift_L11_n_299, B2 => L2_shift_L11_n_204, C => L2_shift_L11_n_295, Z => L2_shift_L11_n_271);
  L2_shift_L11_g12389 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_266, B1 => L2_shift_L11_n_265, ZN => L2_shift_L11_n_270);
  L2_shift_L11_g12390 : OAI221D0BWP7T port map(A1 => L2_shift_L11_n_298, A2 => L2_shift_L11_n_199, B1 => L2_shift_L11_n_209, B2 => L2_shift_L11_n_299, C => L2_shift_L11_n_259, ZN => L2_shift_cell_state_out_shift_pacman(5));
  L2_shift_L11_g12391 : OR3XD1BWP7T port map(A1 => L2_shift_L11_n_292, A2 => L2_shift_L11_n_288, A3 => L2_shift_L11_n_263, Z => L2_shift_L11_n_269);
  L2_shift_L11_g12393 : IAO21D0BWP7T port map(A1 => L2_shift_L11_n_253, A2 => L2_shift_L11_n_306, B => L2_shift_L11_n_293, ZN => L2_shift_L11_n_268);
  L2_shift_L11_g12394 : IAO21D0BWP7T port map(A1 => L2_shift_L11_n_246, A2 => L2_shift_L11_n_305, B => L2_shift_L11_n_292, ZN => L2_shift_L11_n_267);
  L2_shift_L11_g12395 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_298, A2 => L2_shift_L11_n_213, B => L2_shift_L11_n_258, ZN => L2_shift_cell_state_out_shift_pacman(4));
  L2_shift_L11_g12396 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_250, A2 => L2_shift_L11_n_304, B => L2_shift_L11_n_261, ZN => L2_shift_L11_n_266);
  L2_shift_L11_g12397 : CKND1BWP7T port map(I => L2_shift_L11_n_262, ZN => L2_shift_L11_n_263);
  L2_shift_L11_g12398 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_254, A2 => L2_shift_L11_n_302, ZN => L2_shift_L11_n_265);
  L2_shift_L11_g12399 : INR2XD0BWP7T port map(A1 => L2_shift_L11_n_305, B1 => L2_shift_L11_n_245, ZN => L2_shift_L11_n_292);
  L2_shift_L11_g12400 : INR2XD0BWP7T port map(A1 => L2_shift_L11_n_286, B1 => L2_shift_L11_n_247, ZN => L2_shift_L11_n_264);
  L2_shift_L11_g12401 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_251, A2 => L2_shift_L11_n_303, ZN => L2_shift_L11_n_262);
  L2_shift_L11_g12402 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_252, A2 => L2_shift_L11_n_286, ZN => L2_shift_L11_n_289);
  L2_shift_L11_g12403 : INR2XD0BWP7T port map(A1 => L2_shift_L11_n_306, B1 => L2_shift_L11_n_255, ZN => L2_shift_L11_n_293);
  L2_shift_L11_g12405 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_243, A2 => L2_shift_L11_n_210, B1 => L2_shift_L11_n_296, B2 => L2_shift_L11_n_215, ZN => L2_shift_L11_n_259);
  L2_shift_L11_g12406 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_297, A2 => L2_shift_L11_n_217, B => L2_shift_L11_n_258, ZN => L2_shift_cell_state_out_shift_pacman(3));
  L2_shift_L11_g12407 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_249, A2 => L2_shift_L11_n_304, ZN => L2_shift_L11_n_261);
  L2_shift_L11_g12408 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_248, A2 => L2_shift_L11_n_303, ZN => L2_shift_L11_n_288);
  L2_shift_L11_g12409 : INR2XD0BWP7T port map(A1 => L2_shift_L11_n_257, B1 => L2_shift_L11_n_302, ZN => L2_shift_L11_n_287);
  L2_shift_L11_g12410 : CKAN2D1BWP7T port map(A1 => L2_shift_L11_n_244, A2 => L2_county(2), Z => L2_shift_L11_n_290);
  L2_shift_L11_g12411 : OAI22D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_209, B1 => L2_shift_L11_n_405, B2 => L2_shift_L11_n_208, ZN => L2_shift_L11_n_260);
  L2_shift_L11_g12412 : AO22D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_315, B1 => L2_shift_L11_n_314, B2 => L2_shift_L11_n_307, Z => L2_shift_L11_n_257);
  L2_shift_L11_g12413 : AO22D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_311, B1 => L2_shift_L11_n_318, B2 => L2_shift_L11_n_307, Z => L2_shift_L11_n_256);
  L2_shift_L11_g12414 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_321, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_308, ZN => L2_shift_L11_n_255);
  L2_shift_L11_g12415 : AO22D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_314, B1 => L2_shift_L11_n_315, B2 => L2_shift_L11_n_307, Z => L2_shift_L11_n_254);
  L2_shift_L11_g12416 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_308, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_321, ZN => L2_shift_L11_n_253);
  L2_shift_L11_g12417 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_296, B1 => L2_shift_L11_n_230, ZN => L2_shift_L11_n_258);
  L2_shift_L11_g12418 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_307, ZN => L2_shift_L11_n_299);
  L2_shift_L11_g12419 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_307, ZN => L2_shift_L11_n_298);
  L2_shift_L11_g12420 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_317, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_312, ZN => L2_shift_L11_n_252);
  L2_shift_L11_g12421 : AO22D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_313, B1 => L2_shift_L11_n_316, B2 => L2_shift_L11_n_307, Z => L2_shift_L11_n_251);
  L2_shift_L11_g12422 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_310, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_319, ZN => L2_shift_L11_n_250);
  L2_shift_L11_g12423 : AO22D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_319, B1 => L2_shift_L11_n_310, B2 => L2_shift_L11_n_307, Z => L2_shift_L11_n_249);
  L2_shift_L11_g12424 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_316, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_313, ZN => L2_shift_L11_n_248);
  L2_shift_L11_g12425 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_312, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_317, ZN => L2_shift_L11_n_247);
  L2_shift_L11_g12426 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_309, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_320, ZN => L2_shift_L11_n_246);
  L2_shift_L11_g12427 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_320, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_309, ZN => L2_shift_L11_n_245);
  L2_shift_L11_g12428 : AO22D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_318, B1 => L2_shift_L11_n_311, B2 => L2_shift_L11_n_307, Z => L2_shift_L11_n_244);
  L2_shift_L11_g12429 : INVD0BWP7T port map(I => L2_shift_L11_n_297, ZN => L2_shift_L11_n_243);
  L2_shift_L11_g12430 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_307, ZN => L2_shift_L11_n_297);
  L2_shift_L11_g12431 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_307, ZN => L2_shift_L11_n_296);
  L2_shift_L11_g12432 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_241, A2 => L2_shift_L11_n_211, A3 => L2_shift_L11_n_188, A4 => L2_shift_L11_n_223, ZN => L2_shift_L11_n_294);
  L2_shift_L11_g12433 : AOI211XD0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L11_n_228, B => L2_shift_L11_n_242, C => L2_shift_L11_n_231, ZN => L2_shift_L11_n_406);
  L2_shift_L11_g12434 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_218, A2 => L2_shift_L11_n_238, A3 => L2_shift_L11_n_200, A4 => L2_shift_L11_n_224, ZN => L2_shift_L11_n_337);
  L2_shift_L11_g12435 : OR4D1BWP7T port map(A1 => L2_shift_L11_n_202, A2 => L2_shift_L11_n_188, A3 => L2_shift_L11_n_239, A4 => L2_shift_L11_n_211, Z => L2_shift_L11_n_242);
  L2_shift_L11_g12436 : INR4D0BWP7T port map(A1 => L2_shift_L11_n_200, B1 => L2_shift_L11_n_234, B2 => L2_shift_L11_n_240, B3 => L2_shift_L11_n_218, ZN => L2_shift_L11_n_405);
  L2_shift_L11_g12437 : ND3D0BWP7T port map(A1 => L2_shift_L11_n_233, A2 => L2_shift_L11_n_235, A3 => L2_shift_L11_n_202, ZN => L2_shift_L11_n_241);
  L2_shift_L11_g12438 : OAI221D0BWP7T port map(A1 => L2_shift_L11_n_181, A2 => L2_shift_L11_n_220, B1 => L2_shift_L11_n_207, B2 => ycoordinates_int(2), C => L2_shift_L11_n_236, ZN => L2_shift_L11_n_240);
  L2_shift_L11_g12439 : OAI221D0BWP7T port map(A1 => L2_shift_L11_n_172, A2 => L2_shift_L11_n_221, B1 => L2_shift_L11_n_206, B2 => xcoordinates_int(2), C => L2_shift_L11_n_237, ZN => L2_shift_L11_n_239);
  L2_shift_L11_g12440 : OAI221D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_L11_n_225, B1 => L2_shift_L11_n_219, B2 => L2_shift_L11_n_181, C => L2_shift_L11_n_232, ZN => L2_shift_L11_n_238);
  L2_shift_L11_g12441 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_172, A2 => L2_shift_L11_n_221, B1 => xcoordinates_int(2), B2 => L2_shift_L11_n_206, ZN => L2_shift_L11_n_237);
  L2_shift_L11_g12442 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_181, A2 => L2_shift_L11_n_220, B1 => ycoordinates_int(2), B2 => L2_shift_L11_n_207, ZN => L2_shift_L11_n_236);
  L2_shift_L11_g12443 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_171, A2 => L2_shift_L11_n_222, B1 => xcoordinates_int(3), B2 => L2_shift_L11_n_226, ZN => L2_shift_L11_n_235);
  L2_shift_L11_g12444 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_L11_n_229, B1 => ycoordinates_int(3), B2 => L2_shift_L11_n_229, ZN => L2_shift_L11_n_234);
  L2_shift_L11_g12445 : MAOI22D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L11_n_226, B1 => L2_shift_L11_n_171, B2 => L2_shift_L11_n_222, ZN => L2_shift_L11_n_233);
  L2_shift_L11_g12446 : AOI22D0BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_L11_n_225, B1 => L2_shift_L11_n_181, B2 => L2_shift_L11_n_219, ZN => L2_shift_L11_n_232);
  L2_shift_L11_g12447 : NR2D0BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_L11_n_228, ZN => L2_shift_L11_n_231);
  L2_shift_L11_g12448 : OR4D1BWP7T port map(A1 => L2_shift_L11_n_313, A2 => L2_shift_L11_n_314, A3 => L2_shift_L11_n_312, A4 => L2_shift_L11_n_216, Z => L2_shift_L11_n_230);
  L2_shift_L11_g12449 : INVD0BWP7T port map(I => L2_shift_L11_n_307, ZN => L2_shift_L11_n_227);
  L2_shift_L11_g12450 : AOI21D0BWP7T port map(A1 => L2_shift_L11_n_194, A2 => L2_shift_pacman_pos_y(3), B => L2_shift_L11_n_220, ZN => L2_shift_L11_n_229);
  L2_shift_L11_g12451 : AOI21D0BWP7T port map(A1 => L2_shift_L11_n_195, A2 => L2_shift_pacman_pos_x(3), B => L2_shift_L11_n_221, ZN => L2_shift_L11_n_228);
  L2_shift_L11_g12452 : NR3D1BWP7T port map(A1 => L2_shift_L11_n_211, A2 => L2_shift_L11_n_205, A3 => L2_shift_L11_n_171, ZN => L2_shift_L11_n_307);
  L2_shift_L11_g12453 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(2), A2 => L2_shift_L11_n_201, B1 => ycoordinates_int(2), B2 => L2_shift_L11_n_201, ZN => L2_shift_L11_n_224);
  L2_shift_L11_g12454 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(2), A2 => L2_shift_L11_n_198, B1 => xcoordinates_int(2), B2 => L2_shift_L11_n_198, ZN => L2_shift_L11_n_223);
  L2_shift_L11_g12455 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_197, A2 => L2_shift_pacman_pos_x(3), B1 => L2_shift_L11_n_197, B2 => L2_shift_pacman_pos_x(3), ZN => L2_shift_L11_n_226);
  L2_shift_L11_g12456 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_196, A2 => L2_shift_pacman_pos_y(3), B1 => L2_shift_L11_n_196, B2 => L2_shift_pacman_pos_y(3), ZN => L2_shift_L11_n_225);
  L2_shift_L11_g12457 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_197, B1 => L2_shift_pacman_pos_x(3), ZN => L2_shift_L11_n_222);
  L2_shift_L11_g12458 : NR2D0BWP7T port map(A1 => L2_shift_L11_n_195, A2 => L2_shift_pacman_pos_x(3), ZN => L2_shift_L11_n_221);
  L2_shift_L11_g12459 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_194, A2 => L2_shift_pacman_pos_y(3), ZN => L2_shift_L11_n_220);
  L2_shift_L11_g12460 : INR2XD0BWP7T port map(A1 => L2_shift_L11_n_208, B1 => L2_shift_L11_n_210, ZN => L2_shift_L11_n_217);
  L2_shift_L11_g12461 : INR2D1BWP7T port map(A1 => L2_shift_pacman_pos_y(3), B1 => L2_shift_L11_n_196, ZN => L2_shift_L11_n_219);
  L2_shift_L11_g12462 : IND3D1BWP7T port map(A1 => L2_shift_L11_n_205, B1 => L2_shift_L11_n_172, B2 => L2_shift_L11_n_176, ZN => L2_shift_L11_n_218);
  L2_shift_L11_g12463 : INVD1BWP7T port map(I => L2_shift_L11_n_215, ZN => L2_shift_L11_n_216);
  L2_shift_L11_g12464 : INVD0BWP7T port map(I => L2_shift_L11_n_214, ZN => L2_shift_L11_n_213);
  L2_shift_L11_g12465 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_309, A2 => L2_shift_L11_n_311, A3 => L2_shift_L11_n_310, A4 => L2_shift_L11_n_308, ZN => L2_shift_L11_n_215);
  L2_shift_L11_g12466 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_151, A2 => L2_shift_L11_n_191, B => L2_shift_L11_n_199, C => L2_shift_L11_n_192, ZN => L2_shift_L11_n_214);
  L2_shift_L11_g12467 : OA211D0BWP7T port map(A1 => L2_shift_L11_n_150, A2 => L2_shift_L11_n_57, B => L2_shift_L11_n_306, C => L2_shift_L11_n_303, Z => L2_shift_L11_n_212);
  L2_shift_L11_g12468 : IND4D0BWP7T port map(A1 => L2_shift_L11_n_176, B1 => L2_shift_L11_n_181, B2 => L2_shift_L11_n_170, B3 => L2_shift_L11_n_189, ZN => L2_shift_L11_n_211);
  L2_shift_L11_g12469 : OR4D1BWP7T port map(A1 => L2_shift_L11_n_315, A2 => L2_shift_L11_n_318, A3 => L2_shift_L11_n_316, A4 => L2_shift_L11_n_317, Z => L2_shift_L11_n_210);
  L2_shift_L11_g12470 : AO21D0BWP7T port map(A1 => L2_shift_L11_n_193, A2 => L2_shift_L11_n_153, B => L2_shift_L11_n_333, Z => L2_shift_L11_n_204);
  L2_shift_L11_g12471 : AOI211XD0BWP7T port map(A1 => L2_shift_L11_n_185, A2 => L2_shift_L11_n_155, B => L2_shift_L11_n_331, C => L2_shift_L11_n_329, ZN => L2_shift_L11_n_209);
  L2_shift_L11_g12472 : NR3D0BWP7T port map(A1 => L2_shift_L11_n_320, A2 => L2_shift_L11_n_319, A3 => L2_shift_L11_n_321, ZN => L2_shift_L11_n_208);
  L2_shift_L11_g12473 : OA21D0BWP7T port map(A1 => L2_shift_L11_n_164, A2 => L2_shift_L11_n_147, B => L2_shift_L11_n_194, Z => L2_shift_L11_n_207);
  L2_shift_L11_g12474 : OA21D0BWP7T port map(A1 => L2_shift_L11_n_166, A2 => L2_shift_L11_n_148, B => L2_shift_L11_n_195, Z => L2_shift_L11_n_206);
  L2_shift_L11_g12475 : ND4D0BWP7T port map(A1 => L2_shift_L11_n_188, A2 => L2_shift_L11_n_169, A3 => L2_shift_L11_n_142, A4 => L2_shift_L11_n_168, ZN => L2_shift_L11_n_205);
  L2_shift_L11_g12476 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_163, A2 => L2_county(2), B1 => L2_shift_L11_n_163, B2 => L2_county(2), ZN => L2_shift_L11_n_203);
  L2_shift_L11_g12477 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(1), A2 => L2_shift_L11_n_174, B1 => xcoordinates_int(1), B2 => L2_shift_L11_n_174, ZN => L2_shift_L11_n_202);
  L2_shift_L11_g12478 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_156, A2 => L2_shift_pacman_pos_y(2), B1 => L2_shift_L11_n_156, B2 => L2_shift_pacman_pos_y(2), ZN => L2_shift_L11_n_201);
  L2_shift_L11_g12479 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(1), A2 => L2_shift_L11_n_177, B1 => ycoordinates_int(1), B2 => L2_shift_L11_n_177, ZN => L2_shift_L11_n_200);
  L2_shift_L11_g12480 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_193, A2 => L2_shift_L11_n_152, B1 => L2_shift_L11_n_191, B2 => L2_shift_L11_n_154, ZN => L2_shift_L11_n_199);
  L2_shift_L11_g12481 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_157, A2 => L2_shift_pacman_pos_x(2), B1 => L2_shift_L11_n_157, B2 => L2_shift_pacman_pos_x(2), ZN => L2_shift_L11_n_198);
  L2_shift_L11_g12482 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_303, B1 => L2_county(0), ZN => L2_shift_L11_n_302);
  L2_shift_L11_g12483 : OR2D1BWP7T port map(A1 => L2_shift_L11_n_157, A2 => L2_shift_L11_n_148, Z => L2_shift_L11_n_197);
  L2_shift_L11_g12484 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_163, A2 => L2_shift_L11_n_57, ZN => L2_shift_L11_n_304);
  L2_shift_L11_g12485 : OR2D1BWP7T port map(A1 => L2_shift_L11_n_305, A2 => L2_county(0), Z => L2_shift_L11_n_306);
  L2_shift_L11_g12486 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_399, B1 => L2_shift_L11_n_190, ZN => L2_shift_L11_n_295);
  L2_shift_L11_g12487 : OR2D1BWP7T port map(A1 => L2_shift_L11_n_156, A2 => L2_shift_L11_n_147, Z => L2_shift_L11_n_196);
  L2_shift_L11_g12488 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_166, A2 => L2_shift_L11_n_148, ZN => L2_shift_L11_n_195);
  L2_shift_L11_g12489 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_164, A2 => L2_shift_L11_n_147, ZN => L2_shift_L11_n_194);
  L2_shift_L11_g12490 : OAI21D0BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(0), B => L2_county(2), ZN => L2_shift_L11_n_286);
  L2_shift_L11_g12491 : INVD0BWP7T port map(I => L2_shift_L11_n_192, ZN => L2_shift_L11_n_328);
  L2_shift_L11_g12492 : AN2D1BWP7T port map(A1 => L2_shift_L11_n_186, A2 => L2_shift_L11_n_153, Z => L2_shift_L11_n_324);
  L2_shift_L11_g12493 : AN2D1BWP7T port map(A1 => L2_shift_L11_n_185, A2 => L2_shift_L11_state(1), Z => L2_shift_L11_n_330);
  L2_shift_L11_g12494 : AN2D1BWP7T port map(A1 => L2_shift_L11_n_186, A2 => L2_shift_L11_n_152, Z => L2_shift_L11_n_326);
  L2_shift_L11_g12495 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_187, A2 => L2_shift_L11_n_151, ZN => L2_shift_L11_n_322);
  L2_shift_L11_g12496 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_187, A2 => L2_shift_L11_n_154, ZN => L2_shift_L11_n_334);
  L2_shift_L11_g12497 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_187, A2 => L2_shift_L11_n_182, ZN => L2_shift_L11_n_193);
  L2_shift_L11_g12498 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_143, A2 => L2_shift_L11_n_154, ZN => L2_shift_L11_n_331);
  L2_shift_L11_g12499 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_183, A2 => L2_shift_L11_n_153, ZN => L2_shift_L11_n_192);
  L2_shift_L11_g12500 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_184, A2 => L2_shift_L11_n_151, ZN => L2_shift_L11_n_399);
  L2_shift_L11_g12501 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_180, A2 => L2_shift_L11_n_186, ZN => L2_shift_L11_n_191);
  L2_shift_L11_g12502 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_143, A2 => L2_shift_L11_n_151, ZN => L2_shift_L11_n_333);
  L2_shift_L11_g12503 : INR2D1BWP7T port map(A1 => L2_shift_L11_n_186, B1 => L2_shift_L11_n_155, ZN => L2_shift_L11_n_310);
  L2_shift_L11_g12504 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_143, A2 => L2_shift_L11_n_155, ZN => L2_shift_L11_n_317);
  L2_shift_L11_g12505 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_184, A2 => L2_shift_L11_n_162, ZN => L2_shift_L11_n_312);
  L2_shift_L11_g12506 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_184, A2 => L2_shift_L11_n_155, ZN => L2_shift_L11_n_314);
  L2_shift_L11_g12507 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_187, A2 => L2_shift_L11_n_155, ZN => L2_shift_L11_n_320);
  L2_shift_L11_g12508 : AN2D1BWP7T port map(A1 => L2_shift_L11_n_185, A2 => L2_shift_L11_state(4), Z => L2_shift_L11_n_316);
  L2_shift_L11_g12509 : INR2D1BWP7T port map(A1 => L2_shift_L11_n_180, B1 => L2_shift_L11_n_151, ZN => L2_shift_L11_n_327);
  L2_shift_L11_g12510 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_182, A2 => L2_shift_L11_n_151, ZN => L2_shift_L11_n_323);
  L2_shift_L11_g12511 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_182, A2 => L2_shift_L11_n_154, ZN => L2_shift_L11_n_335);
  L2_shift_L11_g12512 : AN2D1BWP7T port map(A1 => L2_shift_L11_n_180, A2 => L2_shift_L11_n_153, Z => L2_shift_L11_n_325);
  L2_shift_L11_g12513 : INR2D1BWP7T port map(A1 => L2_shift_L11_n_185, B1 => L2_shift_L11_n_151, ZN => L2_shift_L11_n_332);
  L2_shift_L11_g12514 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_179, A2 => L2_shift_L11_n_151, ZN => L2_shift_pacman_pos_reset);
  L2_shift_L11_g12515 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_179, A2 => L2_shift_L11_n_154, ZN => L2_shift_L11_n_336);
  L2_shift_L11_g12516 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_152, A2 => L2_shift_L11_n_153, B => L2_shift_L11_n_178, ZN => L2_shift_L11_n_190);
  L2_shift_L11_g12517 : AOI221D0BWP7T port map(A1 => ycoordinates_int(2), A2 => L2_shift_L11_n_147, B1 => L2_shift_L11_n_149, B2 => L2_shift_pacman_pos_y(2), C => L2_shift_L11_n_141, ZN => L2_shift_L11_n_189);
  L2_shift_L11_g12518 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_179, A2 => L2_shift_L11_n_155, ZN => L2_shift_L11_n_329);
  L2_shift_L11_g12519 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_182, A2 => L2_shift_L11_n_155, ZN => L2_shift_L11_n_321);
  L2_shift_L11_g12520 : INR2D1BWP7T port map(A1 => L2_shift_L11_n_180, B1 => L2_shift_L11_n_162, ZN => L2_shift_L11_n_309);
  L2_shift_L11_g12521 : INR2D1BWP7T port map(A1 => L2_shift_L11_n_180, B1 => L2_shift_L11_n_155, ZN => L2_shift_L11_n_311);
  L2_shift_L11_g12522 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_179, A2 => L2_shift_L11_n_162, ZN => L2_shift_L11_n_313);
  L2_shift_L11_g12523 : AN3D1BWP7T port map(A1 => L2_shift_L11_n_161, A2 => L2_shift_L11_state(2), A3 => L2_shift_L11_state(3), Z => L2_shift_L11_n_315);
  L2_shift_L11_g12524 : AN3D1BWP7T port map(A1 => L2_shift_L11_n_161, A2 => L2_shift_L11_state(0), A3 => L2_shift_L11_state(3), Z => L2_shift_L11_n_318);
  L2_shift_L11_g12525 : NR2XD0BWP7T port map(A1 => L2_shift_L11_n_182, A2 => L2_shift_L11_n_162, ZN => L2_shift_L11_n_319);
  L2_shift_L11_g12526 : INVD1BWP7T port map(I => L2_shift_L11_n_183, ZN => L2_shift_L11_n_184);
  L2_shift_L11_g12527 : INVD0BWP7T port map(I => L2_shift_L11_n_179, ZN => L2_shift_L11_n_178);
  L2_shift_L11_g12528 : XNR2D1BWP7T port map(A1 => xcoordinates_int(0), A2 => L2_shift_pacman_pos_x(0), ZN => L2_shift_L11_n_188);
  L2_shift_L11_g12530 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_159, A2 => L2_shift_L11_state(3), ZN => L2_shift_L11_n_187);
  L2_shift_L11_g12531 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_162, A2 => L2_shift_L11_n_158, ZN => L2_shift_L11_n_308);
  L2_shift_L11_g12532 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_158, A2 => L2_shift_L11_state(3), ZN => L2_shift_L11_n_186);
  L2_shift_L11_g12533 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_158, A2 => L2_shift_L11_n_146, ZN => L2_shift_L11_n_185);
  L2_shift_L11_g12534 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_160, A2 => L2_shift_L11_state(3), ZN => L2_shift_L11_n_183);
  L2_shift_L11_g12535 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_165, A2 => L2_shift_L11_state(3), ZN => L2_shift_L11_n_182);
  L2_shift_L11_g12536 : MOAI22D0BWP7T port map(A1 => ycoordinates_int(4), A2 => L2_shift_pacman_pos_y(4), B1 => ycoordinates_int(4), B2 => L2_shift_pacman_pos_y(4), ZN => L2_shift_L11_n_181);
  L2_shift_L11_g12537 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_167, A2 => L2_shift_L11_state(3), ZN => L2_shift_L11_n_180);
  L2_shift_L11_g12538 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_165, A2 => L2_shift_L11_n_146, ZN => L2_shift_L11_n_179);
  L2_shift_L11_g12539 : INVD1BWP7T port map(I => L2_shift_L11_n_172, ZN => L2_shift_L11_n_171);
  L2_shift_L11_g12541 : XNR2D1BWP7T port map(A1 => ycoordinates_int(1), A2 => L2_shift_pacman_pos_y(1), ZN => L2_shift_L11_n_170);
  L2_shift_L11_g12542 : XNR2D1BWP7T port map(A1 => xcoordinates_int(1), A2 => L2_shift_pacman_pos_x(1), ZN => L2_shift_L11_n_169);
  L2_shift_L11_g12543 : MAOI22D0BWP7T port map(A1 => xcoordinates_int(2), A2 => L2_shift_L11_n_148, B1 => xcoordinates_int(2), B2 => L2_shift_L11_n_148, ZN => L2_shift_L11_n_168);
  L2_shift_L11_g12545 : XNR2D1BWP7T port map(A1 => L2_shift_pacman_pos_y(1), A2 => L2_shift_pacman_pos_y(0), ZN => L2_shift_L11_n_177);
  L2_shift_L11_g12546 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(0), A2 => L2_shift_pacman_pos_y(0), Z => L2_shift_L11_n_176);
  L2_shift_L11_g12547 : MOAI22D0BWP7T port map(A1 => L2_shift_L11_n_57, A2 => L2_in_go_y_pos(1), B1 => L2_shift_L11_n_57, B2 => L2_in_go_y_pos(1), ZN => L2_shift_L11_n_175);
  L2_shift_L11_g12548 : CKXOR2D1BWP7T port map(A1 => L2_shift_pacman_pos_x(1), A2 => L2_shift_pacman_pos_x(0), Z => L2_shift_L11_n_174);
  L2_shift_L11_g12549 : MOAI22D0BWP7T port map(A1 => L2_shift_L11_n_150, A2 => L2_in_go_y_pos(1), B1 => L2_shift_L11_n_150, B2 => L2_in_go_y_pos(1), ZN => L2_shift_L11_n_173);
  L2_shift_L11_g12550 : MOAI22D0BWP7T port map(A1 => xcoordinates_int(4), A2 => L2_shift_pacman_pos_x(4), B1 => xcoordinates_int(4), B2 => L2_shift_pacman_pos_x(4), ZN => L2_shift_L11_n_172);
  L2_shift_L11_g12552 : INVD0BWP7T port map(I => L2_shift_L11_n_162, ZN => L2_shift_L11_n_161);
  L2_shift_L11_g12553 : IND2D1BWP7T port map(A1 => L2_shift_L11_state(0), B1 => L2_shift_L11_state(2), ZN => L2_shift_L11_n_167);
  L2_shift_L11_g12554 : NR2XD0BWP7T port map(A1 => L2_shift_pacman_pos_x(1), A2 => L2_shift_pacman_pos_x(0), ZN => L2_shift_L11_n_166);
  L2_shift_L11_g12555 : NR2XD0BWP7T port map(A1 => L2_shift_L11_state(0), A2 => L2_shift_L11_state(2), ZN => L2_shift_L11_n_165);
  L2_shift_L11_g12556 : NR2XD0BWP7T port map(A1 => L2_shift_pacman_pos_y(1), A2 => L2_shift_pacman_pos_y(0), ZN => L2_shift_L11_n_164);
  L2_shift_L11_g12557 : CKND2D1BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(0), ZN => L2_shift_L11_n_163);
  L2_shift_L11_g12558 : ND2D1BWP7T port map(A1 => L2_in_go_y_pos(1), A2 => L2_county(2), ZN => L2_shift_L11_n_303);
  L2_shift_L11_g12559 : ND2D1BWP7T port map(A1 => L2_shift_L11_state(4), A2 => L2_shift_L11_state(1), ZN => L2_shift_L11_n_162);
  L2_shift_L11_g12560 : CKND1BWP7T port map(I => L2_shift_L11_n_159, ZN => L2_shift_L11_n_160);
  L2_shift_L11_g12561 : INVD1BWP7T port map(I => L2_shift_L11_n_154, ZN => L2_shift_L11_n_153);
  L2_shift_L11_g12562 : INVD1BWP7T port map(I => L2_shift_L11_n_152, ZN => L2_shift_L11_n_151);
  L2_shift_L11_g12563 : INR2D1BWP7T port map(A1 => L2_shift_L11_state(0), B1 => L2_shift_L11_state(2), ZN => L2_shift_L11_n_159);
  L2_shift_L11_g12564 : CKND2D1BWP7T port map(A1 => L2_shift_L11_state(0), A2 => L2_shift_L11_state(2), ZN => L2_shift_L11_n_158);
  L2_shift_L11_g12565 : ND2D1BWP7T port map(A1 => L2_shift_pacman_pos_x(1), A2 => L2_shift_pacman_pos_x(0), ZN => L2_shift_L11_n_157);
  L2_shift_L11_g12566 : ND2D1BWP7T port map(A1 => L2_shift_pacman_pos_y(1), A2 => L2_shift_pacman_pos_y(0), ZN => L2_shift_L11_n_156);
  L2_shift_L11_g12568 : IND2D1BWP7T port map(A1 => L2_shift_L11_state(1), B1 => L2_shift_L11_state(4), ZN => L2_shift_L11_n_155);
  L2_shift_L11_g12569 : IND2D1BWP7T port map(A1 => L2_shift_L11_state(4), B1 => L2_shift_L11_state(1), ZN => L2_shift_L11_n_154);
  L2_shift_L11_g12570 : NR2D1BWP7T port map(A1 => L2_shift_L11_state(4), A2 => L2_shift_L11_state(1), ZN => L2_shift_L11_n_152);
  L2_shift_L11_g12574 : INVD0BWP7T port map(I => L2_county(0), ZN => L2_shift_L11_n_150);
  L2_shift_L11_g12575 : INVD0BWP7T port map(I => ycoordinates_int(2), ZN => L2_shift_L11_n_149);
  L2_shift_L11_g12576 : INVD1BWP7T port map(I => L2_shift_pacman_pos_x(2), ZN => L2_shift_L11_n_148);
  L2_shift_L11_g12577 : INVD1BWP7T port map(I => L2_shift_pacman_pos_y(2), ZN => L2_shift_L11_n_147);
  L2_shift_L11_g12581 : INVD1BWP7T port map(I => L2_county(2), ZN => L2_shift_L11_n_57);
  L2_shift_L11_g2 : INR3D0BWP7T port map(A1 => L2_shift_L11_n_268, B1 => L2_shift_L11_n_289, B2 => L2_shift_L11_n_264, ZN => L2_shift_L11_n_144);
  L2_shift_L11_g12582 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_167, B1 => L2_shift_L11_state(3), ZN => L2_shift_L11_n_143);
  L2_shift_L11_g12583 : XNR2D1BWP7T port map(A1 => xcoordinates_int(3), A2 => L2_shift_pacman_pos_x(3), ZN => L2_shift_L11_n_142);
  L2_shift_L11_g12584 : CKXOR2D1BWP7T port map(A1 => ycoordinates_int(3), A2 => L2_shift_pacman_pos_y(3), Z => L2_shift_L11_n_141);
  L2_shift_L11_g12585 : IND2D1BWP7T port map(A1 => L2_in_go_y_pos(1), B1 => L2_shift_L11_n_57, ZN => L2_shift_L11_n_305);
  L2_shift_L11_g10902 : AO211D0BWP7T port map(A1 => L2_pixel_array_to_shift(1), A2 => L2_shift_L11_n_66, B => L2_shift_L11_n_119, C => L2_shift_L11_n_138, Z => L2_shift_pixel_arr_out_shift_pacman(0));
  L2_shift_L11_g10903 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_75, A2 => L2_shift_L11_n_54, B => L2_shift_L11_n_118, C => L2_shift_L11_n_135, ZN => L2_shift_pixel_arr_out_shift_pacman(7));
  L2_shift_L11_g10904 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_74, A2 => L2_shift_L11_n_54, B => L2_shift_L11_n_111, C => L2_shift_L11_n_134, ZN => L2_shift_pixel_arr_out_shift_pacman(6));
  L2_shift_L11_g10905 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_73, A2 => L2_shift_L11_n_54, B => L2_shift_L11_n_137, C => L2_shift_L11_n_116, ZN => L2_shift_pixel_arr_out_shift_pacman(5));
  L2_shift_L11_g10906 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_84, A2 => L2_shift_L11_n_54, B => L2_shift_L11_n_140, C => L2_shift_L11_n_114, ZN => L2_shift_pixel_arr_out_shift_pacman(3));
  L2_shift_L11_g10907 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_70, A2 => L2_shift_L11_n_54, B => L2_shift_L11_n_139, C => L2_shift_L11_n_115, ZN => L2_shift_pixel_arr_out_shift_pacman(4));
  L2_shift_L11_g10908 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_64, A2 => L2_shift_L11_n_54, B => L2_shift_L11_n_136, C => L2_shift_L11_n_113, ZN => L2_shift_pixel_arr_out_shift_pacman(2));
  L2_shift_L11_g10909 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_129, A2 => L2_shift_L11_n_54, B => L2_shift_L11_n_120, C => L2_shift_L11_n_112, ZN => L2_shift_pixel_arr_out_shift_pacman(1));
  L2_shift_L11_g10910 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L11_n_67, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L11_n_66, C => L2_shift_L11_n_133, ZN => L2_shift_L11_n_140);
  L2_shift_L11_g10911 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(4), A2 => L2_shift_L11_n_130, B1 => L2_pixel_array_to_shift(5), B2 => L2_shift_L11_n_66, C => L2_shift_L11_n_103, ZN => L2_shift_L11_n_139);
  L2_shift_L11_g10912 : OAI22D0BWP7T port map(A1 => L2_shift_L11_n_50, A2 => L2_shift_L11_n_132, B1 => L2_shift_L11_n_49, B2 => L2_shift_L11_n_76, ZN => L2_shift_L11_n_138);
  L2_shift_L11_g10913 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L11_n_130, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L11_n_63, C => L2_shift_L11_n_100, ZN => L2_shift_L11_n_137);
  L2_shift_L11_g10914 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(2), A2 => L2_shift_L11_n_130, B1 => L2_pixel_array_to_shift(3), B2 => L2_shift_L11_n_66, C => L2_shift_L11_n_102, ZN => L2_shift_L11_n_136);
  L2_shift_L11_g10915 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L11_n_131, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L11_n_63, ZN => L2_shift_L11_n_135);
  L2_shift_L11_g10916 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(6), A2 => L2_shift_L11_n_130, B1 => L2_pixel_array_to_shift(7), B2 => L2_shift_L11_n_95, ZN => L2_shift_L11_n_134);
  L2_shift_L11_g10917 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L11_n_130, B1 => L2_shift_L11_n_63, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L11_n_133);
  L2_shift_L11_g10918 : AOI221D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_329, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_328, C => L2_shift_L11_n_130, ZN => L2_shift_L11_n_132);
  L2_shift_L11_g10919 : AO221D0BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_322, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_335, C => L2_shift_L11_n_130, Z => L2_shift_L11_n_131);
  L2_shift_L11_g10920 : INVD0BWP7T port map(I => L2_shift_L11_n_130, ZN => L2_shift_L11_n_129);
  L2_shift_L11_g10921 : ND4D0BWP7T port map(A1 => L2_shift_L11_n_128, A2 => L2_shift_L11_n_61, A3 => L2_shift_L11_n_127, A4 => L2_shift_L11_n_407, ZN => L2_shift_L11_n_130);
  L2_shift_L11_g10922 : AOI211XD0BWP7T port map(A1 => L2_shift_L11_n_297, A2 => L2_shift_L11_n_87, B => L2_shift_L11_n_125, C => L2_shift_L11_n_290, ZN => L2_shift_L11_n_128);
  L2_shift_L11_g10923 : AOI211XD0BWP7T port map(A1 => L2_shift_L11_n_296, A2 => L2_shift_L11_n_109, B => L2_shift_L11_n_126, C => L2_shift_L11_n_123, ZN => L2_shift_L11_n_127);
  L2_shift_L11_g10924 : IND4D0BWP7T port map(A1 => L2_shift_L11_n_295, B1 => L2_shift_L11_n_122, B2 => L2_shift_L11_n_81, B3 => L2_shift_L11_n_124, ZN => L2_shift_L11_n_126);
  L2_shift_L11_g10925 : AO211D0BWP7T port map(A1 => L2_shift_L11_n_298, A2 => L2_shift_L11_n_322, B => L2_shift_L11_n_121, C => L2_shift_L11_n_107, Z => L2_shift_L11_n_125);
  L2_shift_L11_g10926 : OAI31D0BWP7T port map(A1 => L2_shift_L11_n_327, A2 => L2_shift_L11_n_328, A3 => L2_shift_L11_n_89, B => L2_shift_L11_n_298, ZN => L2_shift_L11_n_124);
  L2_shift_L11_g10927 : AO211D0BWP7T port map(A1 => L2_shift_L11_n_110, A2 => L2_shift_L11_n_399, B => L2_shift_pacman_pos_reset, C => L2_shift_L11_n_336, Z => L2_shift_shift_clock_reset);
  L2_shift_L11_g10928 : AOI21D0BWP7T port map(A1 => L2_shift_L11_n_88, A2 => L2_shift_L11_n_62, B => L2_shift_L11_n_307, ZN => L2_shift_L11_n_123);
  L2_shift_L11_g10929 : OAI31D0BWP7T port map(A1 => L2_shift_L11_n_335, A2 => L2_shift_L11_n_334, A3 => L2_shift_L11_n_82, B => L2_shift_L11_n_299, ZN => L2_shift_L11_n_122);
  L2_shift_L11_g10930 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_93, B => L2_shift_L11_n_92, ZN => L2_shift_L11_n_121);
  L2_shift_L11_g10931 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L11_n_67, B1 => L2_pixel_array_to_shift(2), B2 => L2_shift_L11_n_66, C => L2_shift_L11_n_108, ZN => L2_shift_L11_n_120);
  L2_shift_L11_g10932 : OAI221D0BWP7T port map(A1 => L2_shift_L11_n_52, A2 => L2_shift_L11_n_86, B1 => L2_shift_L11_n_85, B2 => L2_shift_L11_n_53, C => L2_shift_L11_n_101, ZN => L2_shift_L11_n_119);
  L2_shift_L11_g10933 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L11_n_83, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L11_n_69, C => L2_shift_L11_n_105, ZN => L2_shift_L11_n_118);
  L2_shift_L11_g10935 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L11_n_94, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L11_n_66, ZN => L2_shift_L11_n_116);
  L2_shift_L11_g10936 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L11_n_99, B1 => L2_pixel_array_to_shift(6), B2 => L2_shift_L11_n_67, ZN => L2_shift_L11_n_115);
  L2_shift_L11_g10937 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L11_n_98, B1 => L2_shift_L11_n_49, B2 => L2_shift_L11_n_72, ZN => L2_shift_L11_n_114);
  L2_shift_L11_g10938 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L11_n_96, B1 => L2_shift_L11_n_49, B2 => L2_shift_L11_n_85, ZN => L2_shift_L11_n_113);
  L2_shift_L11_g10939 : MAOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(7), A2 => L2_shift_L11_n_97, B1 => L2_shift_L11_n_49, B2 => L2_shift_L11_n_86, ZN => L2_shift_L11_n_112);
  L2_shift_L11_g10940 : AOI221D0BWP7T port map(A1 => L2_pixel_array_to_shift(5), A2 => L2_shift_L11_n_63, B1 => L2_pixel_array_to_shift(4), B2 => L2_shift_L11_n_83, C => L2_shift_L11_n_104, ZN => L2_shift_L11_n_111);
  L2_shift_L11_g10941 : OR2D1BWP7T port map(A1 => L2_shift_L11_n_403, A2 => L2_shift_L11_n_91, Z => L2_shift_L11_n_110);
  L2_shift_L11_g10942 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => xcoordinates_int(0), Z => L2_shift_pacman_pos_x_new(0));
  L2_shift_L11_g10943 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => xcoordinates_int(3), Z => L2_shift_pacman_pos_x_new(3));
  L2_shift_L11_g10944 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => ycoordinates_int(4), Z => L2_shift_pacman_pos_y_new(4));
  L2_shift_L11_g10945 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => ycoordinates_int(3), Z => L2_shift_pacman_pos_y_new(3));
  L2_shift_L11_g10946 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_311, B1 => L2_shift_L11_n_90, ZN => L2_shift_L11_n_109);
  L2_shift_L11_g10947 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => ycoordinates_int(2), Z => L2_shift_pacman_pos_y_new(2));
  L2_shift_L11_g10948 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => ycoordinates_int(1), Z => L2_shift_pacman_pos_y_new(1));
  L2_shift_L11_g10949 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => xcoordinates_int(4), Z => L2_shift_pacman_pos_x_new(4));
  L2_shift_L11_g10950 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => ycoordinates_int(0), Z => L2_shift_pacman_pos_y_new(0));
  L2_shift_L11_g10951 : OAI22D0BWP7T port map(A1 => L2_shift_L11_n_52, A2 => L2_shift_L11_n_85, B1 => L2_shift_L11_n_53, B2 => L2_shift_L11_n_72, ZN => L2_shift_L11_n_108);
  L2_shift_L11_g10952 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => xcoordinates_int(1), Z => L2_shift_pacman_pos_x_new(1));
  L2_shift_L11_g10953 : AOI21D0BWP7T port map(A1 => L2_shift_L11_n_77, A2 => L2_shift_L11_n_78, B => L2_shift_L11_n_405, ZN => L2_shift_L11_n_107);
  L2_shift_L11_g10954 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_307, A2 => L2_shift_L11_n_79, B => L2_shift_L11_n_80, ZN => L2_shift_L11_n_106);
  L2_shift_L11_g10955 : OAI22D0BWP7T port map(A1 => L2_shift_L11_n_51, A2 => L2_shift_L11_n_73, B1 => L2_shift_L11_n_56, B2 => L2_shift_L11_n_74, ZN => L2_shift_L11_n_105);
  L2_shift_L11_g10956 : AN2D0BWP7T port map(A1 => L2_shift_pacman_pos_load, A2 => xcoordinates_int(2), Z => L2_shift_pacman_pos_x_new(2));
  L2_shift_L11_g10957 : MOAI22D0BWP7T port map(A1 => L2_shift_L11_n_56, A2 => L2_shift_L11_n_73, B1 => L2_pixel_array_to_shift(3), B2 => L2_shift_L11_n_69, ZN => L2_shift_L11_n_104);
  L2_shift_L11_g10958 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L11_n_63, B1 => L2_shift_L11_n_83, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L11_n_103);
  L2_shift_L11_g10959 : OAI22D0BWP7T port map(A1 => L2_shift_L11_n_53, A2 => L2_shift_L11_n_68, B1 => L2_shift_L11_n_52, B2 => L2_shift_L11_n_72, ZN => L2_shift_L11_n_102);
  L2_shift_L11_g10960 : AOI22D0BWP7T port map(A1 => L2_pixel_array_to_shift(2), A2 => L2_shift_L11_n_67, B1 => L2_pixel_array_to_shift(3), B2 => L2_shift_L11_n_71, ZN => L2_shift_L11_n_101);
  L2_shift_L11_g10961 : AO22D0BWP7T port map(A1 => L2_pixel_array_to_shift(3), A2 => L2_shift_L11_n_83, B1 => L2_shift_L11_n_69, B2 => L2_pixel_array_to_shift(2), Z => L2_shift_L11_n_100);
  L2_shift_L11_g10962 : ND2D0BWP7T port map(A1 => L2_shift_L11_n_72, A2 => L2_shift_L11_n_73, ZN => L2_shift_L11_n_99);
  L2_shift_L11_g10963 : ND2D0BWP7T port map(A1 => L2_shift_L11_n_70, A2 => L2_shift_L11_n_85, ZN => L2_shift_L11_n_98);
  L2_shift_L11_g10964 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_64, A2 => L2_shift_L11_n_76, ZN => L2_shift_L11_n_97);
  L2_shift_L11_g10965 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_84, A2 => L2_shift_L11_n_86, ZN => L2_shift_L11_n_96);
  L2_shift_L11_g10966 : ND2D0BWP7T port map(A1 => L2_shift_L11_n_65, A2 => L2_shift_L11_n_75, ZN => L2_shift_L11_n_95);
  L2_shift_L11_g10967 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_68, A2 => L2_shift_L11_n_74, ZN => L2_shift_L11_n_94);
  L2_shift_L11_g10968 : INR2XD0BWP7T port map(A1 => L2_shift_L11_n_399, B1 => L2_shift_L11_n_403, ZN => L2_shift_pacman_pos_load);
  L2_shift_L11_g10969 : AOI222D0BWP7T port map(A1 => L2_shift_L11_n_319, A2 => L2_shift_L11_n_58, B1 => L2_shift_L11_n_321, B2 => L2_shift_L11_n_55, C1 => L2_shift_L11_n_320, C2 => L2_shift_L11_n_59, ZN => L2_shift_L11_n_93);
  L2_shift_L11_g10970 : OAI31D0BWP7T port map(A1 => L2_shift_L11_n_321, A2 => L2_shift_L11_n_320, A3 => L2_shift_L11_n_319, B => L2_shift_L11_n_297, ZN => L2_shift_L11_n_92);
  L2_shift_L11_g10971 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_405, A2 => L2_shift_L11_n_294, A3 => L2_shift_L11_n_406, A4 => L2_shift_L11_n_337, ZN => L2_shift_L11_n_91);
  L2_shift_L11_g10972 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_314, A2 => L2_shift_L11_n_312, A3 => L2_shift_L11_n_310, A4 => L2_shift_L11_n_313, ZN => L2_shift_L11_n_90);
  L2_shift_L11_g10973 : OR4D1BWP7T port map(A1 => L2_shift_L11_n_324, A2 => L2_shift_L11_n_326, A3 => L2_shift_L11_n_323, A4 => L2_shift_L11_n_325, Z => L2_shift_L11_n_89);
  L2_shift_L11_g10974 : AOI222D0BWP7T port map(A1 => L2_shift_L11_n_310, A2 => L2_shift_L11_n_58, B1 => L2_shift_L11_n_314, B2 => L2_shift_L11_n_302, C1 => L2_shift_L11_n_311, C2 => L2_shift_L11_n_57, ZN => L2_shift_L11_n_88);
  L2_shift_L11_g10975 : OR4D1BWP7T port map(A1 => L2_shift_L11_n_318, A2 => L2_shift_L11_n_315, A3 => L2_shift_L11_n_316, A4 => L2_shift_L11_n_317, Z => L2_shift_L11_n_87);
  L2_shift_L11_g10976 : INVD1BWP7T port map(I => L2_shift_L11_n_84, ZN => L2_shift_L11_n_83);
  L2_shift_L11_g10977 : OR3D1BWP7T port map(A1 => L2_shift_L11_n_332, A2 => L2_shift_L11_n_333, A3 => L2_shift_L11_n_331, Z => L2_shift_L11_n_82);
  L2_shift_L11_g10978 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_329, A2 => L2_shift_L11_n_330, B => L2_shift_L11_n_299, ZN => L2_shift_L11_n_81);
  L2_shift_L11_g10979 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_309, A2 => L2_shift_L11_n_308, B => L2_shift_L11_n_296, ZN => L2_shift_L11_n_80);
  L2_shift_L11_g10980 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_55, A2 => L2_shift_L11_n_308, B1 => L2_shift_L11_n_309, B2 => L2_shift_L11_n_59, ZN => L2_shift_L11_n_79);
  L2_shift_L11_g10981 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_318, A2 => L2_shift_L11_n_57, B1 => L2_shift_L11_n_317, B2 => L2_shift_L11_n_286, ZN => L2_shift_L11_n_78);
  L2_shift_L11_g10982 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_302, A2 => L2_shift_L11_n_315, B1 => L2_shift_L11_n_316, B2 => L2_shift_L11_n_303, ZN => L2_shift_L11_n_77);
  L2_shift_L11_g10983 : ND2D1BWP7T port map(A1 => L2_shift_L11_n_60, A2 => cell_type_int(0), ZN => L2_shift_L11_n_403);
  L2_shift_L11_g10984 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_331, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_326, ZN => L2_shift_L11_n_86);
  L2_shift_L11_g10985 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_332, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_325, ZN => L2_shift_L11_n_85);
  L2_shift_L11_g10986 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_327, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_330, ZN => L2_shift_L11_n_84);
  L2_shift_L11_g10987 : INVD0BWP7T port map(I => L2_shift_L11_n_72, ZN => L2_shift_L11_n_71);
  L2_shift_L11_g10988 : INVD1BWP7T port map(I => L2_shift_L11_n_70, ZN => L2_shift_L11_n_69);
  L2_shift_L11_g10989 : INVD1BWP7T port map(I => L2_shift_L11_n_68, ZN => L2_shift_L11_n_67);
  L2_shift_L11_g10990 : INVD1BWP7T port map(I => L2_shift_L11_n_65, ZN => L2_shift_L11_n_66);
  L2_shift_L11_g10991 : INVD1BWP7T port map(I => L2_shift_L11_n_64, ZN => L2_shift_L11_n_63);
  L2_shift_L11_g10992 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_312, A2 => L2_shift_L11_n_286, B1 => L2_shift_L11_n_313, B2 => L2_shift_L11_n_303, ZN => L2_shift_L11_n_62);
  L2_shift_L11_g10993 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_289, A2 => L2_shift_L11_n_293, A3 => L2_shift_L11_n_287, A4 => L2_shift_L11_n_288, ZN => L2_shift_L11_n_61);
  L2_shift_L11_g10994 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_330, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_327, ZN => L2_shift_L11_n_76);
  L2_shift_L11_g10995 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_323, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_334, ZN => L2_shift_L11_n_75);
  L2_shift_L11_g10996 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_324, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_333, ZN => L2_shift_L11_n_74);
  L2_shift_L11_g10997 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_325, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_332, ZN => L2_shift_L11_n_73);
  L2_shift_L11_g10998 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_333, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_324, ZN => L2_shift_L11_n_72);
  L2_shift_L11_g10999 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_326, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_331, ZN => L2_shift_L11_n_70);
  L2_shift_L11_g11000 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_334, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_323, ZN => L2_shift_L11_n_68);
  L2_shift_L11_g11001 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_406, A2 => L2_shift_L11_n_335, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_322, ZN => L2_shift_L11_n_65);
  L2_shift_L11_g11002 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_294, A2 => L2_shift_L11_n_328, B1 => L2_shift_L11_n_307, B2 => L2_shift_L11_n_329, ZN => L2_shift_L11_n_64);
  L2_shift_L11_g11003 : NR2XD0BWP7T port map(A1 => cell_type_int(2), A2 => cell_type_int(1), ZN => L2_shift_L11_n_60);
  L2_shift_L11_g11004 : INVD0BWP7T port map(I => L2_shift_L11_n_305, ZN => L2_shift_L11_n_59);
  L2_shift_L11_g11005 : INVD0BWP7T port map(I => L2_shift_L11_n_304, ZN => L2_shift_L11_n_58);
  L2_shift_L11_g11007 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(2), ZN => L2_shift_L11_n_56);
  L2_shift_L11_g11008 : INVD0BWP7T port map(I => L2_shift_L11_n_306, ZN => L2_shift_L11_n_55);
  L2_shift_L11_g11009 : INVD1BWP7T port map(I => L2_pixel_array_to_shift(1), ZN => L2_shift_L11_n_54);
  L2_shift_L11_g11010 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(4), ZN => L2_shift_L11_n_53);
  L2_shift_L11_g11011 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(5), ZN => L2_shift_L11_n_52);
  L2_shift_L11_g11012 : INVD0BWP7T port map(I => L2_pixel_array_to_shift(3), ZN => L2_shift_L11_n_51);
  L2_shift_L11_g11013 : CKND1BWP7T port map(I => L2_pixel_array_to_shift(7), ZN => L2_shift_L11_n_50);
  L2_shift_L11_g11014 : INVD1BWP7T port map(I => L2_pixel_array_to_shift(6), ZN => L2_shift_L11_n_49);
  L2_shift_L11_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L11_n_48, Q => L2_shift_L11_state(0));
  L2_shift_L11_g10456 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_47, A2 => L2_shift_L11_n_6, A3 => L2_shift_L11_n_15, A4 => L2_shift_L11_n_0, ZN => L2_shift_L11_n_48);
  L2_shift_L11_g10458 : OAI211D1BWP7T port map(A1 => L2_shift_L11_n_2, A2 => L2_shift_L11_n_5, B => L2_shift_L11_n_18, C => L2_shift_L11_n_45, ZN => L2_shift_L11_n_47);
  L2_shift_L11_g10459 : ND4D0BWP7T port map(A1 => L2_shift_L11_n_26, A2 => L2_shift_L11_n_25, A3 => L2_shift_L11_n_41, A4 => L2_shift_L11_n_27, ZN => L2_shift_L11_n_46);
  L2_shift_L11_g10460 : MOAI22D0BWP7T port map(A1 => L2_shift_L11_n_42, A2 => L2_shift_shift_pulse, B1 => L2_shift_L11_n_32, B2 => L2_shift_shift_pulse, ZN => L2_shift_L11_n_45);
  L2_shift_L11_state_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L11_n_43, Q => L2_shift_L11_state(4));
  L2_shift_L11_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L11_n_44, Q => L2_shift_L11_state(1));
  L2_shift_L11_g10463 : IND4D0BWP7T port map(A1 => L2_shift_L11_n_15, B1 => L2_shift_L11_n_12, B2 => L2_shift_L11_n_26, B3 => L2_shift_L11_n_39, ZN => L2_shift_L11_n_44);
  L2_shift_L11_g10464 : IND4D0BWP7T port map(A1 => L2_shift_L11_n_38, B1 => L2_shift_L11_n_16, B2 => L2_shift_L11_n_17, B3 => L2_shift_L11_n_12, ZN => L2_shift_L11_n_43);
  L2_shift_L11_g10465 : IINR4D0BWP7T port map(A1 => L2_shift_L11_n_37, A2 => L2_shift_L11_n_5, B1 => L2_shift_L11_n_399, B2 => L2_shift_L11_n_322, ZN => L2_shift_L11_n_42);
  L2_shift_L11_state_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_shift_L11_n_40, Q => L2_shift_L11_state(2));
  L2_shift_L11_g10467 : AOI221D0BWP7T port map(A1 => L2_shift_L11_n_36, A2 => L2_shift_L11_n_1, B1 => L2_shift_L11_n_322, B2 => L2_shift_L11_n_4, C => L2_shift_L11_n_20, ZN => L2_shift_L11_n_41);
  L2_shift_L11_g10468 : IND4D0BWP7T port map(A1 => L2_shift_L11_n_29, B1 => L2_shift_L11_n_27, B2 => L2_shift_L11_n_31, B3 => L2_shift_L11_n_33, ZN => L2_shift_L11_n_40);
  L2_shift_L11_g10469 : NR3D0BWP7T port map(A1 => L2_shift_L11_n_24, A2 => L2_shift_L11_n_34, A3 => L2_shift_L11_n_29, ZN => L2_shift_L11_n_39);
  L2_shift_L11_g10470 : ND4D0BWP7T port map(A1 => L2_shift_L11_n_30, A2 => L2_shift_L11_n_25, A3 => L2_shift_L11_n_31, A4 => L2_shift_L11_n_19, ZN => L2_shift_L11_n_38);
  L2_shift_L11_g10471 : INR4D0BWP7T port map(A1 => L2_shift_L11_n_32, B1 => L2_shift_L11_n_308, B2 => L2_shift_pacman_pos_reset, B3 => L2_shift_L11_n_336, ZN => L2_shift_L11_n_37);
  L2_shift_L11_g10472 : IND2D1BWP7T port map(A1 => L2_shift_L11_n_334, B1 => L2_shift_L11_n_35, ZN => L2_shift_L11_n_36);
  L2_shift_L11_g10473 : NR4D0BWP7T port map(A1 => L2_shift_L11_n_22, A2 => L2_shift_L11_n_319, A3 => L2_shift_L11_n_320, A4 => L2_shift_L11_n_316, ZN => L2_shift_L11_n_35);
  L2_shift_L11_g10474 : AO221D0BWP7T port map(A1 => L2_shift_L11_n_28, A2 => L2_shift_shift_pulse, B1 => L2_shift_L11_n_23, B2 => L2_shift_L11_n_2, C => L2_shift_L11_n_21, Z => L2_shift_L11_n_34);
  L2_shift_L11_g10475 : AOI222D0BWP7T port map(A1 => L2_shift_L11_n_23, A2 => L2_shift_shift_pulse, B1 => L2_shift_L11_n_8, B2 => L2_shift_L11_n_1, C1 => L2_shift_L11_n_324, C2 => L2_shift_L11_n_4, ZN => L2_shift_L11_n_33);
  L2_shift_L11_g10476 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_28, A2 => L2_shift_L11_n_23, ZN => L2_shift_L11_n_32);
  L2_shift_L11_g10477 : AOI222D0BWP7T port map(A1 => L2_shift_L11_n_11, A2 => L2_shift_L11_n_405, B1 => L2_shift_L11_n_329, B2 => L2_shift_L11_n_4, C1 => L2_shift_L11_n_9, C2 => L2_shift_L11_n_1, ZN => L2_shift_L11_n_30);
  L2_shift_L11_g10478 : AOI211XD0BWP7T port map(A1 => L2_shift_L11_n_311, A2 => L2_shift_L11_n_1, B => L2_shift_L11_n_13, C => L2_shift_L11_n_20, ZN => L2_shift_L11_n_31);
  L2_shift_L11_g10479 : IOA21D1BWP7T port map(A1 => L2_shift_L11_n_325, A2 => L2_shift_L11_n_1, B => L2_shift_L11_n_19, ZN => L2_shift_L11_n_29);
  L2_shift_L11_g10480 : IND3D1BWP7T port map(A1 => L2_shift_L11_n_13, B1 => L2_shift_L11_n_10, B2 => L2_shift_L11_n_17, ZN => L2_shift_L11_n_28);
  L2_shift_L11_g10481 : MAOI22D0BWP7T port map(A1 => L2_shift_L11_n_330, A2 => L2_shift_L11_n_4, B1 => L2_shift_L11_n_14, B2 => L2_shift_L11_n_0, ZN => L2_shift_L11_n_27);
  L2_shift_L11_g10482 : MOAI22D0BWP7T port map(A1 => L2_shift_L11_n_5, A2 => L2_shift_L11_n_3, B1 => L2_shift_L11_n_11, B2 => L2_shift_L11_n_406, ZN => L2_shift_L11_n_24);
  L2_shift_L11_g10483 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_11, A2 => L2_shift_L11_n_294, B1 => L2_shift_L11_n_335, B2 => L2_shift_L11_n_1, ZN => L2_shift_L11_n_26);
  L2_shift_L11_g10484 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_11, A2 => L2_shift_L11_n_337, B1 => L2_shift_L11_n_321, B2 => L2_shift_L11_n_1, ZN => L2_shift_L11_n_25);
  L2_shift_L11_g10485 : AO211D0BWP7T port map(A1 => L2_shift_L11_n_324, A2 => L2_shift_shift_pulse, B => L2_shift_L11_n_323, C => L2_shift_L11_n_318, Z => L2_shift_L11_n_22);
  L2_shift_L11_g10486 : OA21D0BWP7T port map(A1 => L2_shift_L11_n_6, A2 => L2_shift_L11_n_331, B => L2_shift_L11_n_1, Z => L2_shift_L11_n_21);
  L2_shift_L11_g10487 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_7, A2 => L2_shift_L11_n_0, B => L2_shift_L11_n_16, ZN => L2_shift_L11_n_23);
  L2_shift_L11_g10488 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_337, A2 => L2_shift_L11_n_294, B => L2_shift_L11_n_11, ZN => L2_shift_L11_n_18);
  L2_shift_L11_g10489 : AO21D0BWP7T port map(A1 => L2_shift_L11_n_317, A2 => L2_shift_L11_n_1, B => L2_shift_L11_n_15, Z => L2_shift_L11_n_20);
  L2_shift_L11_g10490 : AOI22D0BWP7T port map(A1 => L2_shift_L11_n_308, A2 => L2_shift_L11_n_4, B1 => L2_shift_L11_n_309, B2 => L2_shift_L11_n_1, ZN => L2_shift_L11_n_19);
  L2_shift_L11_g10491 : NR3D0BWP7T port map(A1 => L2_shift_L11_n_331, A2 => L2_shift_L11_n_333, A3 => L2_shift_L11_n_332, ZN => L2_shift_L11_n_14);
  L2_shift_L11_g10492 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_320, A2 => L2_shift_L11_n_314, B => L2_shift_L11_n_1, ZN => L2_shift_L11_n_17);
  L2_shift_L11_g10493 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_312, A2 => L2_shift_L11_n_318, B => L2_shift_L11_n_1, ZN => L2_shift_L11_n_16);
  L2_shift_L11_g10494 : AN2D1BWP7T port map(A1 => L2_shift_L11_n_315, A2 => L2_shift_L11_n_4, Z => L2_shift_L11_n_15);
  L2_shift_L11_g10495 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_326, A2 => L2_shift_L11_n_332, B => L2_shift_L11_n_1, ZN => L2_shift_L11_n_10);
  L2_shift_L11_g10496 : OA21D0BWP7T port map(A1 => L2_shift_L11_n_310, A2 => L2_shift_L11_n_316, B => L2_shift_L11_n_1, Z => L2_shift_L11_n_13);
  L2_shift_L11_g10497 : OAI21D0BWP7T port map(A1 => L2_shift_L11_n_319, A2 => L2_shift_L11_n_313, B => L2_shift_L11_n_1, ZN => L2_shift_L11_n_12);
  L2_shift_L11_g10498 : INR3D0BWP7T port map(A1 => L2_shift_L11_n_399, B1 => L2_shift_L11_n_0, B2 => L2_shift_L11_n_403, ZN => L2_shift_L11_n_11);
  L2_shift_L11_g10499 : AN2D0BWP7T port map(A1 => L2_shift_L11_n_330, A2 => L2_shift_shift_pulse, Z => L2_shift_L11_n_9);
  L2_shift_L11_g10500 : OR2D1BWP7T port map(A1 => L2_shift_L11_n_327, A2 => L2_shift_L11_n_326, Z => L2_shift_L11_n_8);
  L2_shift_L11_g10501 : NR2D0BWP7T port map(A1 => L2_shift_L11_n_328, A2 => L2_shift_L11_n_334, ZN => L2_shift_L11_n_7);
  L2_shift_L11_g10502 : INVD0BWP7T port map(I => L2_shift_L11_n_4, ZN => L2_shift_L11_n_3);
  L2_shift_L11_g10503 : INR2D1BWP7T port map(A1 => L2_shift_L11_n_336, B1 => L2_calc_start_internal, ZN => L2_shift_L11_n_6);
  L2_shift_L11_g10504 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_324, A2 => L2_shift_L11_n_330, ZN => L2_shift_L11_n_5);
  L2_shift_L11_g10505 : NR2D1BWP7T port map(A1 => L2_shift_L11_n_0, A2 => L2_shift_shift_pulse, ZN => L2_shift_L11_n_4);
  L2_shift_L11_g10506 : INVD0BWP7T port map(I => L2_shift_shift_pulse, ZN => L2_shift_L11_n_2);
  L2_shift_L11_drc_bufs10508 : INVD1BWP7T port map(I => L2_shift_L11_n_1, ZN => L2_shift_L11_n_0);
  L2_shift_L11_drc_bufs10509 : INVD0BWP7T port map(I => reset, ZN => L2_shift_L11_n_1);
  L2_shift_L11_state_reg_3 : DFD1BWP7T port map(CP => clk, D => L2_shift_L11_n_46, Q => L2_shift_L11_state(3), QN => L2_shift_L11_n_146);
  L2_shift_L11_g12588 : INR3D0BWP7T port map(A1 => L2_shift_L11_n_261, B1 => L2_shift_L11_n_106, B2 => L2_shift_L11_n_292, ZN => L2_shift_L11_n_407);
  L1_L6b_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L1_L6b_n_5, Q => L1_L6b_state(0));
  L1_L6b_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => L1_L6b_n_4, Q => L1_vc_pulse);
  L1_L6b_g107 : AO211D0BWP7T port map(A1 => L1_L6b_n_2, A2 => L1_L6b_state(0), B => L1_L6b_n_3, C => reset, Z => L1_L6b_n_5);
  L1_L6b_g108 : INR3D0BWP7T port map(A1 => L1_L6b_state(0), B1 => reset, B2 => L1_L6b_n_3, ZN => L1_L6b_n_4);
  L1_L6b_g109 : NR2D0BWP7T port map(A1 => calc_start_game_int, A2 => L1_vc_pulse, ZN => L1_L6b_n_3);
  L1_L6b_g110 : INVD0BWP7T port map(I => calc_start_game_int, ZN => L1_L6b_n_2);
  L1_L3c_IS1_IC1_move_out_reg_2 : LNQD1BWP7T port map(EN => L1_L3c_IS1_IC1_n_34, D => L1_L3c_IS1_IC1_n_23, Q => L1_L3c_move(2));
  L1_L3c_IS1_IC1_g310 : INR2D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_24, B1 => L1_L3c_IS1_IC1_n_25, ZN => L1_L3c_IS1_IC1_n_34);
  L1_L3c_IS1_IC1_g311 : NR3D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_26, A2 => L1_L3c_IS1_IC1_state(2), A3 => L1_L3c_IS1_IC1_state(0), ZN => L1_L3c_IS1_IC1_n_23);
  L1_L3c_IS1_IC1_g312 : ND2D1BWP7T port map(A1 => L1_L3c_IS1_IC1_n_27, A2 => L1_L3c_IS1_IC1_n_26, ZN => L1_L3c_IS1_IC1_n_24);
  L1_L3c_IS1_IC1_g639 : AO21D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_36, A2 => L1_L3c_IS1_IC1_n_15, B => L1_L3c_IS1_IC1_n_19, Z => L1_L3c_IS1_IC1_n_22);
  L1_L3c_IS1_IC1_g640 : AO22D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_36, A2 => L1_L3c_IS1_IC1_n_16, B1 => L1_L3c_IS1_IC1_n_18, B2 => L1_L3c_IS1_IC1_n_1, Z => L1_L3c_IS1_IC1_n_21);
  L1_L3c_IS1_IC1_g641 : AO32D1BWP7T port map(A1 => L1_L3c_IS1_IC1_n_5, A2 => L1_L3c_IS1_IC1_n_17, A3 => L1_L3c_IS1_IC1_n_9, B1 => L1_L3c_IS1_IC1_n_1, B2 => L1_L3c_IS1_IC1_n_8, Z => L1_L3c_IS1_IC1_n_20);
  L1_L3c_IS1_IC1_g642 : NR4D0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3c_IS1_IC1_n_2, A3 => L1_L3c_IS1_IC1_n_12, A4 => L1_L3c_IS1_IC1_n_8, ZN => L1_L3c_IS1_IC1_n_19);
  L1_L3c_IS1_IC1_g643 : INR3D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_9, B1 => L1_L3c_IS1_IC1_n_8, B2 => L1_L3c_IS1_IC1_n_26, ZN => L1_L3c_IS1_IC1_n_18);
  L1_L3c_IS1_IC1_g644 : INVD0BWP7T port map(I => L1_L3c_IS1_IC1_n_16, ZN => L1_L3c_IS1_IC1_n_17);
  L1_L3c_IS1_IC1_g645 : ND2D1BWP7T port map(A1 => L1_L3c_IS1_IC1_n_9, A2 => L1_L3c_IS1_IC1_n_11, ZN => L1_L3c_IS1_IC1_n_15);
  L1_L3c_IS1_IC1_g646 : IND2D1BWP7T port map(A1 => L1_L3c_IS1_IC1_n_12, B1 => L1_L3c_IS1_IC1_n_11, ZN => L1_L3c_IS1_IC1_n_16);
  L1_L3c_IS1_IC1_move_out_reg_0 : LNQD1BWP7T port map(EN => L1_L3c_IS1_IC1_n_34, D => L1_L3c_IS1_IC1_n_7, Q => L1_L3c_move(0));
  L1_L3c_IS1_IC1_move_out_reg_3 : LNQD1BWP7T port map(EN => L1_L3c_IS1_IC1_n_34, D => L1_L3c_IS1_IC1_n_4, Q => L1_L3c_move(3));
  L1_L3c_IS1_IC1_move_out_reg_1 : LNQD1BWP7T port map(EN => L1_L3c_IS1_IC1_n_34, D => L1_L3c_IS1_IC1_n_6, Q => L1_L3c_move(1));
  L1_L3c_IS1_IC1_g652 : INR4D0BWP7T port map(A1 => L1_L3c_IS1_data_intermediate(2), B1 => L1_L3c_IS1_data_intermediate(0), B2 => L1_L3c_IS1_data_intermediate(1), B3 => L1_L3c_IS1_data_intermediate(3), ZN => L1_L3c_IS1_IC1_n_12);
  L1_L3c_IS1_IC1_g653 : IND3D1BWP7T port map(A1 => L1_L3c_IS1_data_intermediate(0), B1 => L1_L3c_IS1_data_intermediate(1), B2 => L1_L3c_IS1_IC1_n_3, ZN => L1_L3c_IS1_IC1_n_11);
  L1_L3c_IS1_IC1_g655 : IND3D1BWP7T port map(A1 => L1_L3c_IS1_data_intermediate(1), B1 => L1_L3c_IS1_data_intermediate(0), B2 => L1_L3c_IS1_IC1_n_3, ZN => L1_L3c_IS1_IC1_n_9);
  L1_L3c_IS1_IC1_g656 : INR4D0BWP7T port map(A1 => L1_L3c_IS1_data_intermediate(3), B1 => L1_L3c_IS1_data_intermediate(0), B2 => L1_L3c_IS1_data_intermediate(1), B3 => L1_L3c_IS1_data_intermediate(2), ZN => L1_L3c_IS1_IC1_n_8);
  L1_L3c_IS1_IC1_g657 : NR2D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_2, A2 => L1_L3c_IS1_IC1_state(1), ZN => L1_L3c_IS1_IC1_n_7);
  L1_L3c_IS1_IC1_g658 : NR2D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_2, A2 => L1_L3c_IS1_IC1_n_26, ZN => L1_L3c_IS1_IC1_n_6);
  L1_L3c_IS1_IC1_g659 : NR3D0BWP7T port map(A1 => L1_L3c_IS1_IC1_n_25, A2 => L1_L3c_IS1_IC1_state(0), A3 => L1_L3c_IS1_IC1_state(1), ZN => L1_L3c_IS1_IC1_n_4);
  L1_L3c_IS1_IC1_g660 : NR3D0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3c_IS1_IC1_n_24, A3 => L1_L3c_IS1_IC1_n_25, ZN => L1_L3c_IS1_IC1_n_5);
  L1_L3c_IS1_IC1_g661 : NR2XD0BWP7T port map(A1 => L1_L3c_IS1_data_intermediate(2), A2 => L1_L3c_IS1_data_intermediate(3), ZN => L1_L3c_IS1_IC1_n_3);
  L1_L3c_IS1_IC1_g663 : ND2D1BWP7T port map(A1 => L1_L3c_IS1_IC1_n_25, A2 => L1_L3c_IS1_IC1_state(0), ZN => L1_L3c_IS1_IC1_n_2);
  L1_L3c_IS1_IC1_g664 : NR2XD0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3c_IS1_IC1_state(2), ZN => L1_L3c_IS1_IC1_n_1);
  L1_L3c_IS1_IC1_state_reg_0 : DFD1BWP7T port map(CP => clk, D => L1_L3c_IS1_IC1_n_22, Q => L1_L3c_IS1_IC1_state(0), QN => L1_L3c_IS1_IC1_n_27);
  L1_L3c_IS1_IC1_state_reg_2 : DFD1BWP7T port map(CP => clk, D => L1_L3c_IS1_IC1_n_20, Q => L1_L3c_IS1_IC1_state(2), QN => L1_L3c_IS1_IC1_n_25);
  L1_L3c_IS1_IC1_state_reg_1 : DFD1BWP7T port map(CP => clk, D => L1_L3c_IS1_IC1_n_21, Q => L1_L3c_IS1_IC1_state(1), QN => L1_L3c_IS1_IC1_n_26);
  L1_L3c_IS1_IC1_g679 : OR2D1BWP7T port map(A1 => L1_L3c_IS1_IC1_n_1, A2 => L1_L3c_IS1_IC1_n_5, Z => L1_L3c_IS1_IC1_n_36);
  L1_L3a_L1_move_out_reg_1 : LNQD1BWP7T port map(EN => L1_L3a_L1_n_34, D => L1_L3a_L1_n_23, Q => L1_L3a_move(1));
  L1_L3a_L1_g310 : NR2D0BWP7T port map(A1 => L1_L3a_L1_n_35, A2 => L1_L3a_L1_n_26, ZN => L1_L3a_L1_n_23);
  L1_L3a_L1_g311 : INR2D0BWP7T port map(A1 => L1_L3a_L1_n_24, B1 => L1_L3a_L1_n_25, ZN => L1_L3a_L1_n_34);
  L1_L3a_L1_g312 : ND2D1BWP7T port map(A1 => L1_L3a_L1_n_25, A2 => L1_L3a_L1_state(0), ZN => L1_L3a_L1_n_35);
  L1_L3a_L1_g313 : ND2D1BWP7T port map(A1 => L1_L3a_L1_n_27, A2 => L1_L3a_L1_n_26, ZN => L1_L3a_L1_n_24);
  L1_L3a_L1_g648 : OR2D1BWP7T port map(A1 => L1_L3a_L1_n_36, A2 => L1_L3a_L1_n_19, Z => L1_L3a_L1_n_22);
  L1_L3a_L1_g649 : AO22D0BWP7T port map(A1 => L1_L3a_L1_n_14, A2 => L1_L3a_L1_n_15, B1 => L1_L3a_L1_n_17, B2 => L1_L3a_L1_n_1, Z => L1_L3a_L1_n_21);
  L1_L3a_L1_g650 : AO32D1BWP7T port map(A1 => L1_L3a_L1_n_7, A2 => L1_L3a_L1_n_16, A3 => L1_L3a_L1_n_10, B1 => L1_L3a_L1_n_1, B2 => L1_L3a_L1_n_9, Z => L1_L3a_L1_n_20);
  L1_L3a_L1_g651 : NR4D0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3a_L1_n_35, A3 => L1_L3a_L1_n_13, A4 => L1_L3a_L1_n_9, ZN => L1_L3a_L1_n_19);
  L1_L3a_L1_g653 : INR3D0BWP7T port map(A1 => L1_L3a_L1_n_10, B1 => L1_L3a_L1_n_9, B2 => L1_L3a_L1_n_26, ZN => L1_L3a_L1_n_17);
  L1_L3a_L1_g654 : INVD0BWP7T port map(I => L1_L3a_L1_n_15, ZN => L1_L3a_L1_n_16);
  L1_L3a_L1_g655 : IND2D1BWP7T port map(A1 => L1_L3a_L1_n_13, B1 => L1_L3a_L1_n_12, ZN => L1_L3a_L1_n_15);
  L1_L3a_L1_move_out_reg_3 : LNQD1BWP7T port map(EN => L1_L3a_L1_n_34, D => L1_L3a_L1_n_5, Q => L1_L3a_move(3));
  L1_L3a_L1_move_out_reg_2 : LNQD1BWP7T port map(EN => L1_L3a_L1_n_34, D => L1_L3a_L1_n_38, Q => L1_L3a_move(2));
  L1_L3a_L1_g659 : INR4D0BWP7T port map(A1 => L1_L3a_data_buffed(2), B1 => L1_L3a_data_buffed(0), B2 => L1_L3a_data_buffed(1), B3 => L1_L3a_data_buffed(3), ZN => L1_L3a_L1_n_13);
  L1_L3a_L1_g660 : IND3D1BWP7T port map(A1 => L1_L3a_data_buffed(0), B1 => L1_L3a_data_buffed(1), B2 => L1_L3a_L1_n_4, ZN => L1_L3a_L1_n_12);
  L1_L3a_L1_g662 : IND3D1BWP7T port map(A1 => L1_L3a_data_buffed(1), B1 => L1_L3a_data_buffed(0), B2 => L1_L3a_L1_n_4, ZN => L1_L3a_L1_n_10);
  L1_L3a_L1_g663 : INR4D0BWP7T port map(A1 => L1_L3a_data_buffed(3), B1 => L1_L3a_data_buffed(0), B2 => L1_L3a_data_buffed(1), B3 => L1_L3a_data_buffed(2), ZN => L1_L3a_L1_n_9);
  L1_L3a_L1_move_out_reg_0 : LNQD1BWP7T port map(EN => L1_L3a_L1_n_34, D => L1_L3a_L1_n_3, Q => L1_L3a_move(0));
  L1_L3a_L1_g667 : NR3D0BWP7T port map(A1 => L1_L3a_L1_n_25, A2 => L1_L3a_L1_state(0), A3 => L1_L3a_L1_state(1), ZN => L1_L3a_L1_n_5);
  L1_L3a_L1_g668 : NR3D0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3a_L1_n_24, A3 => L1_L3a_L1_n_25, ZN => L1_L3a_L1_n_7);
  L1_L3a_L1_g669 : NR2D0BWP7T port map(A1 => L1_L3a_L1_n_35, A2 => L1_L3a_L1_state(1), ZN => L1_L3a_L1_n_3);
  L1_L3a_L1_g670 : NR2XD0BWP7T port map(A1 => L1_L3a_data_buffed(2), A2 => L1_L3a_data_buffed(3), ZN => L1_L3a_L1_n_4);
  L1_L3a_L1_g673 : NR2XD0BWP7T port map(A1 => game_over_out_int, A2 => L1_L3a_L1_state(2), ZN => L1_L3a_L1_n_1);
  L1_L3a_L1_g677 : INVD0BWP7T port map(I => L1_L3a_L1_n_37, ZN => L1_L3a_L1_n_14);
  L1_L3a_L1_g2 : AOI21D0BWP7T port map(A1 => L1_L3a_L1_n_12, A2 => L1_L3a_L1_n_10, B => L1_L3a_L1_n_37, ZN => L1_L3a_L1_n_36);
  L1_L3a_L1_g678 : NR2D1BWP7T port map(A1 => L1_L3a_L1_n_1, A2 => L1_L3a_L1_n_7, ZN => L1_L3a_L1_n_37);
  L1_L3a_L1_state_reg_0 : DFD1BWP7T port map(CP => clk, D => L1_L3a_L1_n_22, Q => L1_L3a_L1_state(0), QN => L1_L3a_L1_n_27);
  L1_L3a_L1_state_reg_2 : DFD1BWP7T port map(CP => clk, D => L1_L3a_L1_n_20, Q => L1_L3a_L1_state(2), QN => L1_L3a_L1_n_25);
  L1_L3a_L1_state_reg_1 : DFD1BWP7T port map(CP => clk, D => L1_L3a_L1_n_21, Q => L1_L3a_L1_state(1), QN => L1_L3a_L1_n_26);
  L1_L3a_L1_g685 : NR3D0BWP7T port map(A1 => L1_L3a_L1_n_26, A2 => L1_L3a_L1_state(0), A3 => L1_L3a_L1_state(2), ZN => L1_L3a_L1_n_38);
  L2_vidcontrol_g2390 : AN2D0BWP7T port map(A1 => L2_vidcontrol_n_60, A2 => L2_vidcontrol_colour_buffer(2), Z => L2_rgb_video(2));
  L2_vidcontrol_g2391 : AN2D0BWP7T port map(A1 => L2_vidcontrol_n_60, A2 => L2_vidcontrol_colour_buffer(1), Z => L2_rgb_video(1));
  L2_vidcontrol_g2392 : AN2D0BWP7T port map(A1 => L2_vidcontrol_n_60, A2 => L2_vidcontrol_colour_buffer(0), Z => L2_rgb_video(0));
  L2_vidcontrol_g2393 : ND4D0BWP7T port map(A1 => L2_vidcontrol_n_59, A2 => L2_vidcontrol_n_56, A3 => L2_vidcontrol_n_58, A4 => L2_vidcontrol_n_57, ZN => L2_vidcontrol_n_60);
  L2_vidcontrol_g2394 : AO21D0BWP7T port map(A1 => L2_vidcontrol_n_54, A2 => L2_vidcontrol_n_55, B => L2_vidcontrol_n_52, Z => L2_reset_current_block_vertical);
  L2_vidcontrol_g2395 : INR3D0BWP7T port map(A1 => L2_vidcontrol_n_54, B1 => L2_vidcontrol_n_41, B2 => L2_vidcontrol_n_55, ZN => L2_en_current_block_vertical);
  L2_vidcontrol_g2396 : OR2D0BWP7T port map(A1 => L2_vidcontrol_n_54, A2 => L2_vidcontrol_n_52, Z => L2_reset_county_video);
  L2_vidcontrol_g2397 : NR3D0BWP7T port map(A1 => L2_vidcontrol_n_53, A2 => L2_vidcontrol_n_45, A3 => L2_vidcontrol_n_41, ZN => L2_en_county_video);
  L2_vidcontrol_g2398 : AOI22D0BWP7T port map(A1 => L2_vidcontrol_n_82, A2 => L2_vidcontrol_pixel_arr_buffer(7), B1 => L2_vidcontrol_n_79, B2 => L2_vidcontrol_pixel_arr_buffer(5), ZN => L2_vidcontrol_n_59);
  L2_vidcontrol_g2399 : AOI22D0BWP7T port map(A1 => L2_vidcontrol_n_76, A2 => L2_vidcontrol_pixel_arr_buffer(1), B1 => L2_vidcontrol_n_11, B2 => L2_vidcontrol_pixel_arr_buffer(3), ZN => L2_vidcontrol_n_58);
  L2_vidcontrol_g2400 : AOI22D0BWP7T port map(A1 => L2_en_current_block_horizontal_video, A2 => L2_vidcontrol_pixel_arr_buffer(6), B1 => L2_vidcontrol_n_78, B2 => L2_vidcontrol_pixel_arr_buffer(4), ZN => L2_vidcontrol_n_57);
  L2_vidcontrol_g2401 : AOI22D0BWP7T port map(A1 => L2_vidcontrol_n_3, A2 => L2_vidcontrol_pixel_arr_buffer(0), B1 => L2_vidcontrol_n_77, B2 => L2_vidcontrol_pixel_arr_buffer(2), ZN => L2_vidcontrol_n_56);
  L2_vidcontrol_g2402 : OR2D0BWP7T port map(A1 => L2_vidcontrol_n_52, A2 => L2_vidcontrol_n_47, Z => L2_reset_current_block_horizontal_video);
  L2_vidcontrol_g2403 : INR2XD0BWP7T port map(A1 => L2_current_block_vertical(3), B1 => L2_vidcontrol_n_52, ZN => ycoordinates_int(3));
  L2_vidcontrol_g2404 : INR2XD0BWP7T port map(A1 => L2_current_block_vertical(2), B1 => L2_vidcontrol_n_52, ZN => ycoordinates_int(2));
  L2_vidcontrol_g2405 : INR2XD0BWP7T port map(A1 => L2_current_block_vertical(1), B1 => L2_vidcontrol_n_52, ZN => ycoordinates_int(1));
  L2_vidcontrol_g2406 : INR2XD0BWP7T port map(A1 => L2_current_block_vertical(0), B1 => L2_vidcontrol_n_52, ZN => ycoordinates_int(0));
  L2_vidcontrol_g2407 : ND2D0BWP7T port map(A1 => L2_vidcontrol_n_51, A2 => L2_vidcontrol_n_53, ZN => L2_reset_dual_pixel_y_video);
  L2_vidcontrol_g2408 : INR2D1BWP7T port map(A1 => L2_current_block_vertical(4), B1 => L2_vidcontrol_n_52, ZN => ycoordinates_int(4));
  L2_vidcontrol_g2409 : AN2D1BWP7T port map(A1 => L2_vidcontrol_n_51, A2 => L2_current_block_horizontal(2), Z => xcoordinates_int(2));
  L2_vidcontrol_g2410 : INR3D0BWP7T port map(A1 => L2_vidcontrol_n_47, B1 => L2_dual_pixel_y, B2 => L2_vidcontrol_n_41, ZN => L2_en_dual_pixel_y_video);
  L2_vidcontrol_g2411 : AN2D1BWP7T port map(A1 => L2_vidcontrol_n_51, A2 => L2_current_block_horizontal(4), Z => xcoordinates_int(4));
  L2_vidcontrol_g2412 : AN2D1BWP7T port map(A1 => L2_vidcontrol_n_51, A2 => L2_current_block_horizontal(3), Z => xcoordinates_int(3));
  L2_vidcontrol_g2413 : AN2D1BWP7T port map(A1 => L2_vidcontrol_n_51, A2 => L2_current_block_horizontal(0), Z => xcoordinates_int(0));
  L2_vidcontrol_g2414 : CKAN2D1BWP7T port map(A1 => L2_vidcontrol_n_51, A2 => L2_current_block_horizontal(1), Z => xcoordinates_int(1));
  L2_vidcontrol_g2415 : INR2D1BWP7T port map(A1 => L2_current_block_vertical(4), B1 => L2_vidcontrol_n_50, ZN => L2_vidcontrol_n_55);
  L2_vidcontrol_g2416 : INR2XD0BWP7T port map(A1 => L2_vidcontrol_n_45, B1 => L2_vidcontrol_n_53, ZN => L2_vidcontrol_n_54);
  L2_vidcontrol_g2417 : NR2D1BWP7T port map(A1 => L2_vidcontrol_n_49, A2 => L2_vidcontrol_state(1), ZN => L2_vidcontrol_n_78);
  L2_vidcontrol_g2418 : INR2D1BWP7T port map(A1 => L2_vidcontrol_state(1), B1 => L2_vidcontrol_n_46, ZN => L2_vidcontrol_n_11);
  L2_vidcontrol_g2419 : INR2D1BWP7T port map(A1 => L2_vidcontrol_state(1), B1 => L2_vidcontrol_n_49, ZN => L2_vidcontrol_n_77);
  L2_vidcontrol_g2420 : ND2D1BWP7T port map(A1 => L2_vidcontrol_n_47, A2 => L2_dual_pixel_y, ZN => L2_vidcontrol_n_53);
  L2_vidcontrol_g2421 : INVD1BWP7T port map(I => L2_vidcontrol_n_52, ZN => L2_vidcontrol_n_51);
  L2_vidcontrol_g2422 : AOI31D0BWP7T port map(A1 => L2_current_block_vertical(2), A2 => L2_current_block_vertical(1), A3 => L2_current_block_vertical(0), B => L2_current_block_vertical(3), ZN => L2_vidcontrol_n_50);
  L2_vidcontrol_g2423 : NR3D0BWP7T port map(A1 => L2_vidcontrol_n_42, A2 => L2_vidcontrol_n_39, A3 => L2_vidcontrol_state(2), ZN => L2_vidcontrol_n_82);
  L2_vidcontrol_g2424 : NR3D0BWP7T port map(A1 => L2_vidcontrol_n_43, A2 => L2_vidcontrol_n_39, A3 => L2_vidcontrol_state(2), ZN => L2_en_current_block_horizontal_video);
  L2_vidcontrol_g2425 : NR2D1BWP7T port map(A1 => L2_vidcontrol_n_46, A2 => L2_vidcontrol_state(1), ZN => L2_vidcontrol_n_79);
  L2_vidcontrol_g2426 : OR2D1BWP7T port map(A1 => L2_vidcontrol_n_123, A2 => L2_vidcontrol_n_72, Z => L2_vidcontrol_n_52);
  L2_vidcontrol_g2427 : INVD0BWP7T port map(I => L2_vidcontrol_n_3, ZN => L2_vidcontrol_n_124);
  L2_vidcontrol_g2428 : NR2XD0BWP7T port map(A1 => L2_vidcontrol_n_41, A2 => L2_vidcontrol_state(3), ZN => L2_vidcontrol_n_83);
  L2_vidcontrol_g2429 : IND2D1BWP7T port map(A1 => L2_vidcontrol_n_43, B1 => L2_vidcontrol_state(2), ZN => L2_vidcontrol_n_49);
  L2_vidcontrol_g2430 : NR2D1BWP7T port map(A1 => L2_vidcontrol_n_41, A2 => L2_vidcontrol_n_44, ZN => L2_vidcontrol_n_3);
  L2_vidcontrol_g2431 : NR2XD0BWP7T port map(A1 => L2_vidcontrol_n_125, A2 => L2_vidcontrol_n_44, ZN => L2_vidcontrol_n_47);
  L2_vidcontrol_g2432 : NR2XD0BWP7T port map(A1 => L2_vidcontrol_n_41, A2 => L2_vidcontrol_n_42, ZN => L2_vidcontrol_n_123);
  L2_vidcontrol_g2433 : CKAN2D1BWP7T port map(A1 => L2_vidcontrol_n_41, A2 => L2_vidcontrol_state(3), Z => L2_vidcontrol_n_72);
  L2_vidcontrol_g2434 : IND2D1BWP7T port map(A1 => L2_vidcontrol_n_42, B1 => L2_vidcontrol_state(2), ZN => L2_vidcontrol_n_46);
  L2_vidcontrol_g2435 : AN3D1BWP7T port map(A1 => L2_county(0), A2 => L2_county(2), A3 => L2_in_go_y_pos(1), Z => L2_vidcontrol_n_45);
  L2_vidcontrol_g2436 : NR3D0BWP7T port map(A1 => L2_vidcontrol_n_41, A2 => L2_vidcontrol_n_40, A3 => L2_vidcontrol_state(0), ZN => L2_vidcontrol_n_76);
  L2_vidcontrol_g2437 : ND2D1BWP7T port map(A1 => L2_current_block_horizontal(3), A2 => L2_current_block_horizontal(4), ZN => L2_vidcontrol_n_125);
  L2_vidcontrol_g2438 : ND2D1BWP7T port map(A1 => L2_vidcontrol_state(0), A2 => L2_vidcontrol_state(3), ZN => L2_vidcontrol_n_44);
  L2_vidcontrol_g2439 : ND2D1BWP7T port map(A1 => L2_vidcontrol_n_40, A2 => L2_vidcontrol_state(0), ZN => L2_vidcontrol_n_43);
  L2_vidcontrol_g2440 : IND2D1BWP7T port map(A1 => L2_vidcontrol_state(0), B1 => L2_vidcontrol_n_40, ZN => L2_vidcontrol_n_42);
  L2_vidcontrol_g2441 : IND2D1BWP7T port map(A1 => L2_vidcontrol_state(2), B1 => L2_vidcontrol_n_39, ZN => L2_vidcontrol_n_41);
  L2_vidcontrol_colour_buffer_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_37, Q => L2_vidcontrol_colour_buffer(0));
  L2_vidcontrol_colour_buffer_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_38, Q => L2_vidcontrol_colour_buffer(1));
  L2_vidcontrol_colour_buffer_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_36, Q => L2_vidcontrol_colour_buffer(2));
  L2_vidcontrol_pixel_arr_buffer_reg_6 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_32, Q => L2_vidcontrol_pixel_arr_buffer(6));
  L2_vidcontrol_pixel_arr_buffer_reg_5 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_34, Q => L2_vidcontrol_pixel_arr_buffer(5));
  L2_vidcontrol_pixel_arr_buffer_reg_4 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_33, Q => L2_vidcontrol_pixel_arr_buffer(4));
  L2_vidcontrol_pixel_arr_buffer_reg_7 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_31, Q => L2_vidcontrol_pixel_arr_buffer(7));
  L2_vidcontrol_g2122 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_29, A2 => L2_vidcontrol_colour_buffer(1), B1 => L2_vidcontrol_n_28, B2 => L2_sprite_colour(1), Z => L2_vidcontrol_n_38);
  L2_vidcontrol_g2124 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_29, A2 => L2_vidcontrol_colour_buffer(0), B1 => L2_vidcontrol_n_28, B2 => L2_sprite_colour(0), Z => L2_vidcontrol_n_37);
  L2_vidcontrol_g2125 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_29, A2 => L2_vidcontrol_colour_buffer(2), B1 => L2_vidcontrol_n_28, B2 => L2_sprite_colour(2), Z => L2_vidcontrol_n_36);
  L2_vidcontrol_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_30, Q => L2_vidcontrol_state(0));
  L2_vidcontrol_state_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => L2_vidcontrol_n_19, D => L2_vidcontrol_n_21, Q => L2_vidcontrol_state(2));
  L2_vidcontrol_pixel_arr_buffer_reg_3 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_26, Q => L2_vidcontrol_pixel_arr_buffer(3));
  L2_vidcontrol_pixel_arr_buffer_reg_0 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_23, Q => L2_vidcontrol_pixel_arr_buffer(0));
  L2_vidcontrol_pixel_arr_buffer_reg_1 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_24, Q => L2_vidcontrol_pixel_arr_buffer(1));
  L2_vidcontrol_pixel_arr_buffer_reg_2 : DFQD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_25, Q => L2_vidcontrol_pixel_arr_buffer(2));
  L2_vidcontrol_g2133 : OAI21D0BWP7T port map(A1 => L2_vidcontrol_n_16, A2 => L2_vidcontrol_n_5, B => L2_vidcontrol_n_27, ZN => L2_vidcontrol_n_35);
  L2_vidcontrol_g2134 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_126, A2 => L2_vidcontrol_pixel_arr_buffer(5), B1 => L2_vidcontrol_n_18, B2 => L2_pixel_array_shifted(5), Z => L2_vidcontrol_n_34);
  L2_vidcontrol_g2135 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_126, A2 => L2_vidcontrol_pixel_arr_buffer(4), B1 => L2_vidcontrol_n_18, B2 => L2_pixel_array_shifted(4), Z => L2_vidcontrol_n_33);
  L2_vidcontrol_g2136 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_126, A2 => L2_vidcontrol_pixel_arr_buffer(6), B1 => L2_vidcontrol_n_18, B2 => L2_pixel_array_shifted(6), Z => L2_vidcontrol_n_32);
  L2_vidcontrol_g2137 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_126, A2 => L2_vidcontrol_pixel_arr_buffer(7), B1 => L2_vidcontrol_n_18, B2 => L2_pixel_array_shifted(7), Z => L2_vidcontrol_n_31);
  L2_vidcontrol_g2138 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_21, A2 => L2_vidcontrol_n_20, B1 => L2_vidcontrol_n_4, B2 => L2_vidcontrol_n_15, Z => L2_vidcontrol_n_30);
  L2_vidcontrol_g2139 : OAI21D0BWP7T port map(A1 => L2_vidcontrol_n_8, A2 => L2_vidcontrol_n_82, B => L2_vidcontrol_n_21, ZN => L2_vidcontrol_n_27);
  L2_vidcontrol_g2140 : INR2D1BWP7T port map(A1 => L2_vidcontrol_n_22, B1 => reset, ZN => L2_vidcontrol_n_29);
  L2_vidcontrol_g2141 : NR2D1BWP7T port map(A1 => L2_vidcontrol_n_22, A2 => reset, ZN => L2_vidcontrol_n_28);
  L2_vidcontrol_g2142 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_14, A2 => L2_vidcontrol_pixel_arr_buffer(3), B1 => L2_vidcontrol_n_12, B2 => L2_pixel_array_shifted(3), Z => L2_vidcontrol_n_26);
  L2_vidcontrol_g2143 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_14, A2 => L2_vidcontrol_pixel_arr_buffer(2), B1 => L2_vidcontrol_n_12, B2 => L2_pixel_array_shifted(2), Z => L2_vidcontrol_n_25);
  L2_vidcontrol_g2144 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_14, A2 => L2_vidcontrol_pixel_arr_buffer(1), B1 => L2_vidcontrol_n_12, B2 => L2_pixel_array_shifted(1), Z => L2_vidcontrol_n_24);
  L2_vidcontrol_g2145 : AO22D0BWP7T port map(A1 => L2_vidcontrol_n_14, A2 => L2_vidcontrol_pixel_arr_buffer(0), B1 => L2_vidcontrol_n_12, B2 => L2_pixel_array_shifted(0), Z => L2_vidcontrol_n_23);
  L2_vidcontrol_g2146 : NR4D0BWP7T port map(A1 => L2_en_current_block_horizontal_video, A2 => L2_vidcontrol_n_77, A3 => L2_vidcontrol_n_78, A4 => L2_vidcontrol_n_72, ZN => L2_vidcontrol_n_20);
  L2_vidcontrol_g2147 : OR3D1BWP7T port map(A1 => L2_vidcontrol_n_79, A2 => L2_en_current_block_horizontal_video, A3 => L2_vidcontrol_n_8, Z => L2_vidcontrol_n_19);
  L2_vidcontrol_g2148 : NR2XD0BWP7T port map(A1 => L2_vidcontrol_n_13, A2 => L2_vidcontrol_n_123, ZN => L2_vidcontrol_n_22);
  L2_vidcontrol_g2149 : NR2XD0BWP7T port map(A1 => L2_vidcontrol_n_5, A2 => L2_vidcontrol_n_13, ZN => L2_vidcontrol_n_21);
  L2_vidcontrol_g2150 : AOI22D0BWP7T port map(A1 => L2_n_536, A2 => L2_vidcontrol_n_6, B1 => L2_vidcontrol_n_3, B2 => L2_vidcontrol_n_125, ZN => L2_vidcontrol_n_16);
  L2_vidcontrol_g2151 : OAI22D0BWP7T port map(A1 => L2_n_536, A2 => L2_vidcontrol_n_7, B1 => L2_vidcontrol_n_124, B2 => L2_vidcontrol_n_125, ZN => L2_vidcontrol_n_15);
  L2_vidcontrol_g2152 : IAO21D0BWP7T port map(A1 => L2_vidcontrol_n_11, A2 => L2_vidcontrol_n_83, B => reset, ZN => L2_vidcontrol_n_18);
  L2_vidcontrol_g2154 : INR2D1BWP7T port map(A1 => L2_vidcontrol_n_10, B1 => reset, ZN => L2_vidcontrol_n_14);
  L2_vidcontrol_g2155 : ND2D1BWP7T port map(A1 => L2_vidcontrol_n_7, A2 => L2_vidcontrol_n_124, ZN => L2_vidcontrol_n_13);
  L2_vidcontrol_g2156 : NR2XD0BWP7T port map(A1 => L2_vidcontrol_n_10, A2 => reset, ZN => L2_vidcontrol_n_12);
  L2_vidcontrol_g2157 : OR2D1BWP7T port map(A1 => L2_vidcontrol_n_76, A2 => L2_vidcontrol_n_77, Z => L2_vidcontrol_n_9);
  L2_vidcontrol_g2159 : NR2XD0BWP7T port map(A1 => L2_vidcontrol_n_82, A2 => L2_vidcontrol_n_83, ZN => L2_vidcontrol_n_10);
  L2_vidcontrol_g2160 : INVD0BWP7T port map(I => L2_vidcontrol_n_7, ZN => L2_vidcontrol_n_6);
  L2_vidcontrol_g2161 : INVD0BWP7T port map(I => L2_vidcontrol_n_4, ZN => L2_vidcontrol_n_5);
  L2_vidcontrol_g2162 : OR2D1BWP7T port map(A1 => L2_vidcontrol_n_11, A2 => L2_vidcontrol_n_78, Z => L2_vidcontrol_n_8);
  L2_vidcontrol_g2163 : ND2D1BWP7T port map(A1 => L2_vidcontrol_n_83, A2 => L2_vidcontrol_state(0), ZN => L2_vidcontrol_n_7);
  L2_vidcontrol_g2164 : NR2XD0BWP7T port map(A1 => L2_user_reset_new, A2 => reset, ZN => L2_vidcontrol_n_4);
  L2_vidcontrol_g2 : NR3D0BWP7T port map(A1 => L2_vidcontrol_n_83, A2 => L2_vidcontrol_n_11, A3 => reset, ZN => L2_vidcontrol_n_126);
  L2_vidcontrol_state_reg_3 : DFKCND1BWP7T port map(CP => clk, CN => L2_vidcontrol_n_9, D => L2_vidcontrol_n_21, Q => L2_vidcontrol_state(3), QN => L2_vidcontrol_n_40);
  L2_vidcontrol_state_reg_1 : DFD1BWP7T port map(CP => clk, D => L2_vidcontrol_n_35, Q => L2_vidcontrol_state(1), QN => L2_vidcontrol_n_39);
  L1_L3c_IS1_IB1_FF1_data_out_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_pacman(3), D => L1_L3c_IS1_IB1_FF1_n_0, Q => L1_L3c_IS1_IB1_data_intermediate(3));
  L1_L3c_IS1_IB1_FF1_data_out_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_pacman(2), D => L1_L3c_IS1_IB1_FF1_n_0, Q => L1_L3c_IS1_IB1_data_intermediate(2));
  L1_L3c_IS1_IB1_FF1_data_out_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_pacman(0), D => L1_L3c_IS1_IB1_FF1_n_0, Q => L1_L3c_IS1_IB1_data_intermediate(0));
  L1_L3c_IS1_IB1_FF1_data_out_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => dir_pacman(1), D => L1_L3c_IS1_IB1_FF1_n_0, Q => L1_L3c_IS1_IB1_data_intermediate(1));
  L1_L3c_IS1_IB1_FF1_g7 : INVD1BWP7T port map(I => game_over_out_int, ZN => L1_L3c_IS1_IB1_FF1_n_0);
  L1_L3c_IS1_IB1_FF2_data_out_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3c_IS1_IB1_data_intermediate(3), D => L1_L3c_IS1_IB1_FF2_n_0, Q => L1_L3c_IS1_data_intermediate(3));
  L1_L3c_IS1_IB1_FF2_data_out_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3c_IS1_IB1_data_intermediate(2), D => L1_L3c_IS1_IB1_FF2_n_0, Q => L1_L3c_IS1_data_intermediate(2));
  L1_L3c_IS1_IB1_FF2_data_out_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3c_IS1_IB1_data_intermediate(0), D => L1_L3c_IS1_IB1_FF2_n_0, Q => L1_L3c_IS1_data_intermediate(0));
  L1_L3c_IS1_IB1_FF2_data_out_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => L1_L3c_IS1_IB1_data_intermediate(1), D => L1_L3c_IS1_IB1_FF2_n_0, Q => L1_L3c_IS1_data_intermediate(1));
  L1_L3c_IS1_IB1_FF2_g7 : INVD1BWP7T port map(I => game_over_out_int, ZN => L1_L3c_IS1_IB1_FF2_n_0);

end synthesised;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity d_flipflop_1bit is
  	port ( 	
		clk		: in std_logic;
		signal_in 	: in std_logic;
	        signal_out 	: out std_logic
	);
end entity d_flipflop_1bit;



configuration shift_control_behaviour_cfg of shift_control is
   for behaviour
   end for;
end shift_control_behaviour_cfg;

library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of score_control is
begin
end behaviour;


configuration pacman_position_reg_behavioural_cfg of pacman_position_reg is
   for behavioural
   end for;
end pacman_position_reg_behavioural_cfg;

configuration score_counter_behaviour_cfg of score_counter is
   for behaviour
   end for;
end score_counter_behaviour_cfg;

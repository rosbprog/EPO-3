library IEEE;
use IEEE.std_logic_1164.ALL;

entity total_system_tb is
end total_system_tb;


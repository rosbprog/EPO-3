configuration pacman_cont_behaviour_cfg of pacman_cont is
   for behaviour
   end for;
end pacman_cont_behaviour_cfg;

configuration plus_one_behaviour_cfg of plus_one is
   for behaviour
   end for;
end plus_one_behaviour_cfg;

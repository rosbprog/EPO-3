configuration score_sprite_behavioural_cfg of score_sprite is
   for behavioural
   end for;
end score_sprite_behavioural_cfg;

configuration new_counter_behaviour_cfg of new_counter is
   for behaviour
   end for;
end new_counter_behaviour_cfg;
